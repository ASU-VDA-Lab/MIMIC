module fake_netlist_6_121_n_1152 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1152);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1152;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_1119;
wire n_344;
wire n_946;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_1075;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_72),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_181),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_68),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_16),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_24),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_21),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_131),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_134),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_91),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_32),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_151),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_109),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_169),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_139),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_120),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_157),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_88),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_6),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_105),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_86),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_128),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_144),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_93),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_74),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_83),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_54),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_115),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_116),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_92),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_164),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_45),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_36),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_80),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_155),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_70),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_133),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_226),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_228),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_229),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_268),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_260),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_244),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_262),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_277),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_243),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_256),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_287),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_256),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_240),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_222),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_224),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_225),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_249),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_230),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_255),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_231),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_248),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_232),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_276),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_318),
.B1(n_295),
.B2(n_302),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_313),
.Y(n_346)
);

OAI22x1_ASAP7_75t_R g347 ( 
.A1(n_319),
.A2(n_266),
.B1(n_281),
.B2(n_252),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

NOR2x1_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_223),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g351 ( 
.A(n_332),
.B(n_264),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_324),
.A2(n_286),
.B1(n_289),
.B2(n_290),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_233),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_308),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_234),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_309),
.B(n_0),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_323),
.B(n_0),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_325),
.B(n_285),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_292),
.B(n_248),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_294),
.B(n_235),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_329),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_329),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_292),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_1),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_236),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_297),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_304),
.A2(n_316),
.B(n_315),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_331),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_237),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_324),
.A2(n_283),
.B1(n_280),
.B2(n_275),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_241),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_293),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_340),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_293),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_393),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_338),
.B1(n_340),
.B2(n_302),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_395),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_305),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_305),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_356),
.B(n_311),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_372),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_248),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_394),
.B(n_311),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_346),
.B(n_242),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_371),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_SL g415 ( 
.A(n_388),
.B(n_245),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_342),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_301),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_371),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_369),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_368),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_394),
.B(n_246),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_361),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

NOR2x1p5_ASAP7_75t_L g429 ( 
.A(n_374),
.B(n_247),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_341),
.B(n_250),
.Y(n_430)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_379),
.A2(n_322),
.B(n_301),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_353),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_355),
.B(n_257),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_384),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_390),
.Y(n_445)
);

BUFx6f_ASAP7_75t_SL g446 ( 
.A(n_351),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_353),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

OR2x2_ASAP7_75t_SL g449 ( 
.A(n_357),
.B(n_322),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_343),
.B(n_259),
.C(n_258),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_274),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_385),
.B(n_270),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_369),
.B(n_271),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_392),
.B(n_2),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_365),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_348),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_351),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

NOR2x1p5_ASAP7_75t_L g467 ( 
.A(n_375),
.B(n_358),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_349),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_359),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_448),
.Y(n_470)
);

INVx4_ASAP7_75t_SL g471 ( 
.A(n_442),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_387),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_392),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_453),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_424),
.B(n_350),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_370),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_387),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_444),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_413),
.B(n_360),
.Y(n_484)
);

OR2x2_ASAP7_75t_SL g485 ( 
.A(n_450),
.B(n_368),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_363),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

XNOR2x2_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_367),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_430),
.B(n_2),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_408),
.B(n_33),
.Y(n_493)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_3),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_455),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_408),
.B(n_34),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_416),
.B(n_35),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_359),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_443),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_432),
.B(n_3),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_4),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_414),
.B(n_37),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_447),
.B(n_366),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_415),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_415),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_454),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_426),
.B(n_38),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_464),
.B(n_364),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_469),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_370),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_454),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_423),
.B(n_364),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_409),
.A2(n_370),
.B(n_376),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_446),
.B(n_366),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_4),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_431),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_414),
.B(n_40),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_398),
.B(n_42),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_402),
.B(n_406),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_421),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_421),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_43),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_423),
.B(n_5),
.Y(n_547)
);

XOR2x2_ASAP7_75t_L g548 ( 
.A(n_445),
.B(n_410),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_423),
.B(n_452),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_400),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_452),
.B(n_5),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_420),
.B(n_376),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_420),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_490),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_509),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_452),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_481),
.B(n_472),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_521),
.A2(n_446),
.B1(n_467),
.B2(n_425),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_499),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_500),
.B(n_411),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_492),
.A2(n_457),
.B1(n_446),
.B2(n_409),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_492),
.A2(n_456),
.B1(n_463),
.B2(n_460),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_485),
.A2(n_449),
.B1(n_433),
.B2(n_429),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_482),
.A2(n_456),
.B1(n_463),
.B2(n_460),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_411),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_501),
.B(n_400),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_473),
.B(n_521),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_495),
.B(n_400),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_549),
.B(n_459),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_474),
.B(n_439),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_470),
.B(n_459),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_516),
.B(n_439),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_530),
.B(n_401),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_516),
.A2(n_401),
.B1(n_403),
.B2(n_428),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_529),
.A2(n_439),
.B(n_403),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_496),
.B(n_401),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_403),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_489),
.B(n_428),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_542),
.B(n_428),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_436),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_507),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_518),
.B(n_439),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_479),
.A2(n_436),
.B1(n_427),
.B2(n_407),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_479),
.A2(n_436),
.B1(n_427),
.B2(n_407),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_407),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_478),
.B(n_407),
.Y(n_593)
);

O2A1O1Ixp5_ASAP7_75t_L g594 ( 
.A1(n_480),
.A2(n_466),
.B(n_437),
.C(n_427),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_504),
.B(n_407),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_483),
.B(n_427),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_486),
.B(n_427),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_538),
.B(n_437),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_517),
.B(n_437),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_538),
.B(n_466),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_511),
.B(n_6),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_498),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_476),
.B(n_7),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_491),
.A2(n_466),
.B1(n_9),
.B2(n_10),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_487),
.B(n_8),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_8),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_511),
.B(n_10),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_488),
.B(n_11),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_532),
.B(n_11),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_529),
.B(n_44),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_510),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_515),
.B(n_12),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_484),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_536),
.B(n_520),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_484),
.B(n_12),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_536),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_539),
.B(n_13),
.Y(n_620)
);

BUFx8_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_540),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_471),
.B(n_46),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_582),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_531),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_571),
.B(n_548),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_569),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_561),
.B(n_614),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_603),
.A2(n_541),
.B1(n_546),
.B2(n_494),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_563),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_601),
.B(n_543),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_560),
.B(n_503),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_556),
.B(n_471),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_588),
.B(n_567),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_599),
.Y(n_639)
);

AO22x1_ASAP7_75t_L g640 ( 
.A1(n_605),
.A2(n_493),
.B1(n_502),
.B2(n_523),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_577),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_604),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_595),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_559),
.B(n_471),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_544),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_577),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_583),
.B(n_545),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_575),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_575),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_609),
.B(n_551),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_577),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_617),
.B(n_552),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_573),
.B(n_554),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_621),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_512),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_577),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_611),
.B(n_513),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_588),
.B(n_514),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_562),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_601),
.B(n_550),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_587),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_570),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_572),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_612),
.A2(n_533),
.B(n_535),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_584),
.B(n_522),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_558),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_608),
.B(n_526),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_565),
.B(n_533),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_581),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_593),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_622),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_610),
.B(n_527),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_622),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_568),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_576),
.B(n_537),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_686),
.A2(n_612),
.B(n_566),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_659),
.A2(n_620),
.A3(n_602),
.B(n_600),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_670),
.B(n_597),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_679),
.A2(n_623),
.B(n_579),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_630),
.A2(n_578),
.B1(n_606),
.B2(n_591),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_624),
.B(n_601),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_667),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_667),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_659),
.A2(n_598),
.A3(n_579),
.B(n_594),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_672),
.A2(n_590),
.B(n_574),
.Y(n_697)
);

NOR2x1_ASAP7_75t_SL g698 ( 
.A(n_641),
.B(n_622),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_643),
.Y(n_699)
);

AOI211x1_ASAP7_75t_L g700 ( 
.A1(n_637),
.A2(n_619),
.B(n_15),
.C(n_16),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_647),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_633),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_L g703 ( 
.A1(n_635),
.A2(n_14),
.B(n_17),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_629),
.A2(n_525),
.B(n_48),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_675),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_658),
.B(n_525),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_679),
.A2(n_670),
.B(n_637),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_651),
.A2(n_49),
.B(n_47),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_648),
.A2(n_674),
.B(n_661),
.Y(n_709)
);

OAI22x1_ASAP7_75t_L g710 ( 
.A1(n_665),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_710)
);

AOI21x1_ASAP7_75t_SL g711 ( 
.A1(n_654),
.A2(n_18),
.B(n_19),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_635),
.A2(n_20),
.B(n_21),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_629),
.A2(n_127),
.B(n_220),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_657),
.A2(n_125),
.B(n_219),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_636),
.A2(n_124),
.B(n_218),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_632),
.B(n_22),
.C(n_23),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_657),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_675),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_638),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_639),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_641),
.A2(n_130),
.B(n_217),
.Y(n_721)
);

OAI22x1_ASAP7_75t_L g722 ( 
.A1(n_628),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_641),
.A2(n_129),
.B(n_216),
.Y(n_723)
);

OA22x2_ASAP7_75t_L g724 ( 
.A1(n_677),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_724)
);

AOI21xp33_ASAP7_75t_L g725 ( 
.A1(n_632),
.A2(n_29),
.B(n_30),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_658),
.Y(n_726)
);

NAND2x1p5_ASAP7_75t_L g727 ( 
.A(n_624),
.B(n_50),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_669),
.A2(n_135),
.B(n_215),
.Y(n_728)
);

OAI21x1_ASAP7_75t_SL g729 ( 
.A1(n_683),
.A2(n_132),
.B(n_214),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_647),
.B(n_51),
.Y(n_730)
);

BUFx12f_ASAP7_75t_L g731 ( 
.A(n_658),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_642),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_653),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_676),
.B(n_29),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_641),
.A2(n_136),
.B(n_52),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_676),
.B(n_30),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_626),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_683),
.B(n_625),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_625),
.B(n_53),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_684),
.A2(n_671),
.B(n_681),
.C(n_663),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_645),
.B(n_55),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_631),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_678),
.A2(n_56),
.B(n_57),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_687),
.A2(n_58),
.B(n_59),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_678),
.A2(n_60),
.B(n_61),
.Y(n_746)
);

NAND2x1_ASAP7_75t_L g747 ( 
.A(n_673),
.B(n_62),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_63),
.B(n_64),
.Y(n_748)
);

OAI21x1_ASAP7_75t_SL g749 ( 
.A1(n_698),
.A2(n_655),
.B(n_650),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_716),
.A2(n_685),
.B1(n_634),
.B2(n_646),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_690),
.B(n_685),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_699),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_690),
.B(n_685),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_682),
.B(n_680),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_735),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_717),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_704),
.A2(n_673),
.B(n_680),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_730),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_688),
.A2(n_634),
.B(n_666),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_726),
.B(n_656),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_702),
.Y(n_761)
);

OAI22x1_ASAP7_75t_L g762 ( 
.A1(n_716),
.A2(n_646),
.B1(n_650),
.B2(n_649),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_703),
.A2(n_634),
.B(n_666),
.C(n_626),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_730),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_SL g765 ( 
.A(n_708),
.B(n_664),
.C(n_640),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_738),
.B(n_725),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_724),
.A2(n_685),
.B1(n_666),
.B2(n_656),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_712),
.A2(n_668),
.B1(n_627),
.B2(n_660),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_735),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_707),
.A2(n_668),
.B(n_644),
.C(n_660),
.Y(n_770)
);

AO32x2_ASAP7_75t_L g771 ( 
.A1(n_719),
.A2(n_664),
.A3(n_660),
.B1(n_652),
.B2(n_647),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_691),
.A2(n_660),
.B(n_652),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_744),
.A2(n_652),
.B(n_647),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_713),
.A2(n_652),
.B(n_644),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_731),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_693),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_745),
.A2(n_627),
.B(n_66),
.C(n_67),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_698),
.A2(n_65),
.A3(n_69),
.B(n_71),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_741),
.A2(n_627),
.B(n_75),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_714),
.A2(n_627),
.B(n_76),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_743),
.B(n_73),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_717),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_693),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_720),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_739),
.B(n_77),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_697),
.A2(n_78),
.B(n_79),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_728),
.A2(n_221),
.B(n_82),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_692),
.A2(n_212),
.B(n_87),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_742),
.A2(n_81),
.B(n_89),
.C(n_90),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_732),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_746),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_791)
);

NOR2x1_ASAP7_75t_SL g792 ( 
.A(n_706),
.B(n_97),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_733),
.Y(n_793)
);

BUFx12f_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_694),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_695),
.B(n_98),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_740),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_715),
.A2(n_711),
.B(n_748),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_721),
.A2(n_103),
.A3(n_104),
.B(n_106),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_723),
.A2(n_211),
.B(n_108),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_729),
.A2(n_107),
.B(n_110),
.C(n_111),
.Y(n_802)
);

OA21x2_ASAP7_75t_L g803 ( 
.A1(n_736),
.A2(n_718),
.B(n_705),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_747),
.A2(n_113),
.B(n_114),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_730),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_701),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_701),
.A2(n_117),
.B(n_118),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_700),
.B(n_119),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_689),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_689),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_701),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_727),
.Y(n_812)
);

O2A1O1Ixp5_ASAP7_75t_SL g813 ( 
.A1(n_700),
.A2(n_121),
.B(n_122),
.C(n_123),
.Y(n_813)
);

AO31x2_ASAP7_75t_L g814 ( 
.A1(n_689),
.A2(n_137),
.A3(n_138),
.B(n_140),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_696),
.A2(n_209),
.B(n_142),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_696),
.A2(n_141),
.B(n_143),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_734),
.A2(n_145),
.B(n_147),
.C(n_148),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_696),
.A2(n_149),
.B(n_150),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_737),
.B(n_152),
.C(n_153),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_710),
.A2(n_154),
.B(n_156),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_793),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_784),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_760),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_765),
.A2(n_722),
.B1(n_159),
.B2(n_160),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_758),
.A2(n_158),
.B1(n_161),
.B2(n_163),
.Y(n_825)
);

INVx6_ASAP7_75t_L g826 ( 
.A(n_794),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_766),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_820),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_761),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_SL g830 ( 
.A1(n_758),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_SL g831 ( 
.A1(n_758),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_776),
.B(n_182),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_775),
.Y(n_833)
);

HB1xp67_ASAP7_75t_SL g834 ( 
.A(n_752),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_790),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_809),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_767),
.B(n_186),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_796),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_755),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_769),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_764),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_803),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_756),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_783),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_763),
.B(n_754),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_811),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_782),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_806),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_810),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_764),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_806),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_764),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_814),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_771),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_803),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_812),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_795),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_805),
.Y(n_858)
);

INVx3_ASAP7_75t_SL g859 ( 
.A(n_751),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_SL g860 ( 
.A1(n_787),
.A2(n_195),
.B1(n_199),
.B2(n_200),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_750),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_753),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_749),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_770),
.A2(n_204),
.B1(n_777),
.B2(n_768),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_819),
.A2(n_788),
.B1(n_792),
.B2(n_808),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_781),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_785),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_814),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_762),
.Y(n_869)
);

INVx6_ASAP7_75t_L g870 ( 
.A(n_797),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_757),
.Y(n_871)
);

BUFx5_ASAP7_75t_L g872 ( 
.A(n_786),
.Y(n_872)
);

INVx4_ASAP7_75t_SL g873 ( 
.A(n_778),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_771),
.Y(n_874)
);

BUFx4_ASAP7_75t_R g875 ( 
.A(n_771),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_774),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_773),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_817),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_816),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_759),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_772),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_798),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_807),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_778),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_836),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_874),
.B(n_778),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_835),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_839),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_879),
.A2(n_818),
.B(n_815),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_856),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_836),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_840),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_849),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_853),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_853),
.A2(n_799),
.B(n_779),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_868),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_842),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_845),
.A2(n_780),
.B(n_801),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_855),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_838),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_880),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_822),
.B(n_813),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_877),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_843),
.B(n_800),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_871),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_847),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_821),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_884),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_876),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_876),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_865),
.A2(n_789),
.B(n_791),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_876),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_875),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_846),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_864),
.A2(n_804),
.B(n_802),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_873),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_852),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_869),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_854),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_834),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_873),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_854),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_872),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_SL g925 ( 
.A1(n_878),
.A2(n_800),
.B1(n_867),
.B2(n_883),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_881),
.B(n_863),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_829),
.B(n_881),
.Y(n_927)
);

BUFx4f_ASAP7_75t_SL g928 ( 
.A(n_833),
.Y(n_928)
);

HB1xp67_ASAP7_75t_SL g929 ( 
.A(n_848),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_882),
.A2(n_878),
.B1(n_824),
.B2(n_860),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_872),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_823),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_870),
.B(n_844),
.Y(n_933)
);

BUFx5_ASAP7_75t_L g934 ( 
.A(n_872),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_858),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_906),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_885),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_885),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_911),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_891),
.Y(n_940)
);

AO21x2_ASAP7_75t_L g941 ( 
.A1(n_889),
.A2(n_837),
.B(n_861),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_887),
.B(n_859),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_911),
.B(n_832),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_886),
.B(n_872),
.Y(n_944)
);

AO21x2_ASAP7_75t_L g945 ( 
.A1(n_889),
.A2(n_825),
.B(n_841),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_891),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_895),
.A2(n_872),
.B(n_828),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_890),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_893),
.Y(n_949)
);

NAND2x1_ASAP7_75t_L g950 ( 
.A(n_926),
.B(n_862),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_899),
.A2(n_827),
.B(n_862),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_906),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_893),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_894),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_894),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_921),
.B(n_857),
.Y(n_957)
);

AO21x1_ASAP7_75t_SL g958 ( 
.A1(n_922),
.A2(n_923),
.B(n_920),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_924),
.B(n_826),
.Y(n_960)
);

AO21x2_ASAP7_75t_L g961 ( 
.A1(n_897),
.A2(n_866),
.B(n_830),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_900),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_897),
.A2(n_866),
.B(n_831),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_886),
.B(n_850),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_900),
.B(n_826),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_888),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_902),
.B(n_870),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_930),
.A2(n_851),
.B1(n_912),
.B2(n_925),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_902),
.B(n_907),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_917),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_898),
.B(n_904),
.Y(n_971)
);

AO21x2_ASAP7_75t_L g972 ( 
.A1(n_931),
.A2(n_896),
.B(n_909),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_950),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_948),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_944),
.B(n_914),
.Y(n_975)
);

AO31x2_ASAP7_75t_L g976 ( 
.A1(n_959),
.A2(n_922),
.A3(n_917),
.B(n_931),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_944),
.B(n_914),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_948),
.Y(n_978)
);

AND2x4_ASAP7_75t_SL g979 ( 
.A(n_960),
.B(n_926),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_955),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_944),
.B(n_923),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_955),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_955),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_956),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_965),
.B(n_915),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_956),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_956),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_959),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_936),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_970),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_953),
.B(n_913),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_970),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_962),
.B(n_898),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_953),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_936),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_936),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_952),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_952),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_985),
.B(n_942),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_975),
.B(n_965),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_983),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_975),
.B(n_965),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_977),
.B(n_960),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_988),
.Y(n_1005)
);

INVx5_ASAP7_75t_SL g1006 ( 
.A(n_991),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_977),
.B(n_942),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_981),
.B(n_967),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_981),
.B(n_990),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_988),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_993),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_993),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_980),
.A2(n_967),
.B(n_972),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_990),
.B(n_960),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_978),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_992),
.B(n_960),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1007),
.B(n_997),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1005),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1013),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1013),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1000),
.A2(n_968),
.B1(n_961),
.B2(n_963),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_1008),
.B(n_973),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_1015),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1010),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1004),
.B(n_973),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1004),
.B(n_973),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_L g1027 ( 
.A(n_1015),
.B(n_919),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_1002),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_1009),
.B(n_979),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1018),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_1014),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_1001),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_1027),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_950),
.Y(n_1034)
);

NOR2x1p5_ASAP7_75t_L g1035 ( 
.A(n_1022),
.B(n_935),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1024),
.B(n_1001),
.Y(n_1036)
);

NAND2x1_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_1009),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_1037),
.B(n_932),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_R g1039 ( 
.A(n_1032),
.B(n_932),
.Y(n_1039)
);

AO221x2_ASAP7_75t_L g1040 ( 
.A1(n_1030),
.A2(n_1020),
.B1(n_1019),
.B2(n_929),
.C(n_1021),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_1029),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1031),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_1021),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1035),
.A2(n_968),
.B1(n_1026),
.B2(n_1017),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1043),
.B(n_1036),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1042),
.B(n_1011),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1041),
.B(n_1034),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_SL g1048 ( 
.A1(n_1039),
.A2(n_957),
.B(n_933),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1040),
.B(n_1012),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1038),
.B(n_1003),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_1043),
.A2(n_1020),
.B1(n_1019),
.B2(n_1028),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1042),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1053),
.A2(n_1028),
.B1(n_1015),
.B2(n_964),
.C(n_992),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_1006),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1049),
.B(n_1055),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1046),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1050),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1045),
.B(n_1014),
.Y(n_1063)
);

OAI322xp33_ASAP7_75t_L g1064 ( 
.A1(n_1053),
.A2(n_974),
.A3(n_927),
.B1(n_1002),
.B2(n_964),
.C1(n_1016),
.C2(n_918),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1061),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1061),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1059),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1057),
.B(n_935),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1058),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1062),
.B(n_1048),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1060),
.B(n_1052),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1065),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1066),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1067),
.Y(n_1075)
);

AOI322xp5_ASAP7_75t_L g1076 ( 
.A1(n_1070),
.A2(n_1056),
.A3(n_1063),
.B1(n_1064),
.B2(n_964),
.C1(n_1016),
.C2(n_974),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1072),
.B(n_1069),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1074),
.B(n_1071),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1073),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1076),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1072),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1078),
.B(n_928),
.Y(n_1083)
);

NOR3x1_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_927),
.C(n_951),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1079),
.B(n_978),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1077),
.B(n_890),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1081),
.A2(n_960),
.B1(n_1006),
.B2(n_948),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1080),
.A2(n_1006),
.B1(n_961),
.B2(n_963),
.Y(n_1088)
);

NAND4xp25_ASAP7_75t_L g1089 ( 
.A(n_1087),
.B(n_943),
.C(n_910),
.D(n_913),
.Y(n_1089)
);

OAI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_1083),
.A2(n_979),
.B(n_926),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1085),
.B(n_916),
.C(n_899),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1086),
.B(n_991),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1088),
.B(n_916),
.C(n_951),
.Y(n_1093)
);

OA211x2_ASAP7_75t_L g1094 ( 
.A1(n_1090),
.A2(n_1084),
.B(n_958),
.C(n_969),
.Y(n_1094)
);

NAND4xp25_ASAP7_75t_L g1095 ( 
.A(n_1089),
.B(n_943),
.C(n_910),
.D(n_969),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_961),
.B(n_963),
.C(n_945),
.Y(n_1096)
);

NAND5xp2_ASAP7_75t_L g1097 ( 
.A(n_1093),
.B(n_905),
.C(n_903),
.D(n_961),
.E(n_963),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_1091),
.B(n_951),
.C(n_908),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1090),
.B(n_958),
.C(n_998),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1092),
.B(n_994),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1090),
.A2(n_991),
.B1(n_998),
.B2(n_999),
.C(n_945),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_926),
.B(n_991),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_945),
.B(n_947),
.C(n_941),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_1095),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1101),
.A2(n_999),
.B1(n_994),
.B2(n_995),
.C(n_989),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_1097),
.B(n_994),
.Y(n_1106)
);

NOR3x2_ASAP7_75t_L g1107 ( 
.A(n_1094),
.B(n_947),
.C(n_945),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1098),
.B(n_1096),
.C(n_982),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1099),
.B(n_941),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_1099),
.B(n_994),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_1108),
.B(n_982),
.C(n_986),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_1104),
.B(n_939),
.C(n_905),
.Y(n_1112)
);

NAND4xp75_ASAP7_75t_L g1113 ( 
.A(n_1106),
.B(n_980),
.C(n_987),
.D(n_986),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1109),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1110),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_L g1116 ( 
.A(n_1102),
.B(n_947),
.Y(n_1116)
);

AOI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1107),
.A2(n_996),
.B1(n_995),
.B2(n_989),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1105),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1103),
.Y(n_1119)
);

NAND4xp25_ASAP7_75t_L g1120 ( 
.A(n_1104),
.B(n_943),
.C(n_903),
.D(n_939),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1104),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_SL g1122 ( 
.A(n_1104),
.B(n_987),
.C(n_996),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_943),
.Y(n_1123)
);

AOI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1115),
.A2(n_966),
.B(n_984),
.C(n_983),
.Y(n_1124)
);

AOI22x1_ASAP7_75t_L g1125 ( 
.A1(n_1119),
.A2(n_984),
.B1(n_939),
.B2(n_966),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_SL g1126 ( 
.A(n_1114),
.B(n_901),
.C(n_949),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1118),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1113),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1111),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1117),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1127),
.A2(n_1122),
.B1(n_1112),
.B2(n_1120),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_939),
.B2(n_947),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1129),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1128),
.A2(n_937),
.B1(n_949),
.B2(n_946),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1130),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1125),
.A2(n_953),
.B1(n_937),
.B2(n_938),
.Y(n_1136)
);

OAI22x1_ASAP7_75t_L g1137 ( 
.A1(n_1131),
.A2(n_1126),
.B1(n_1124),
.B2(n_953),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1133),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1138),
.A2(n_1132),
.B(n_1136),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1140),
.Y(n_1141)
);

AOI21xp33_ASAP7_75t_SL g1142 ( 
.A1(n_1141),
.A2(n_1139),
.B(n_1137),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_1134),
.B1(n_940),
.B2(n_954),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_946),
.B1(n_954),
.B2(n_940),
.Y(n_1144)
);

AO22x2_ASAP7_75t_L g1145 ( 
.A1(n_1143),
.A2(n_938),
.B1(n_962),
.B2(n_952),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_941),
.B1(n_934),
.B2(n_972),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_941),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1146),
.B(n_896),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_SL g1149 ( 
.A1(n_1145),
.A2(n_901),
.B(n_892),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1147),
.B(n_976),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_1148),
.B1(n_1149),
.B2(n_888),
.C(n_892),
.Y(n_1151)
);

AOI211xp5_ASAP7_75t_L g1152 ( 
.A1(n_1151),
.A2(n_971),
.B(n_962),
.C(n_904),
.Y(n_1152)
);


endmodule