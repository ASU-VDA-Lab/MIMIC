module fake_jpeg_18827_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_23),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_42),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_70),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_43),
.B1(n_35),
.B2(n_42),
.Y(n_63)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_63),
.B(n_98),
.CI(n_26),
.CON(n_132),
.SN(n_132)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_34),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_78),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_18),
.B1(n_41),
.B2(n_33),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_18),
.B1(n_41),
.B2(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_36),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_33),
.B1(n_39),
.B2(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_39),
.B1(n_22),
.B2(n_17),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_95),
.B1(n_52),
.B2(n_26),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_89),
.Y(n_130)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_27),
.B1(n_17),
.B2(n_29),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_100),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_99),
.B(n_101),
.C(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_21),
.B1(n_31),
.B2(n_28),
.Y(n_93)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_26),
.A3(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_21),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2x1p5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_46),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_122),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_28),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_112),
.C(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_23),
.C(n_49),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_126),
.B(n_129),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_26),
.A3(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_77),
.B1(n_84),
.B2(n_97),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_68),
.A2(n_26),
.B(n_23),
.C(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_90),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_99),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_142),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_23),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_144),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_68),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_76),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_97),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_143),
.B(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_78),
.B1(n_82),
.B2(n_63),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_154),
.B1(n_83),
.B2(n_91),
.Y(n_172)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_151),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_116),
.B(n_131),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_162),
.B(n_87),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_63),
.C(n_79),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_100),
.C(n_87),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_62),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_90),
.B1(n_74),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_155),
.B1(n_141),
.B2(n_133),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_109),
.A2(n_93),
.B1(n_67),
.B2(n_80),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_107),
.A2(n_103),
.B1(n_131),
.B2(n_123),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_102),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_122),
.B(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_89),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_8),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_164),
.B(n_6),
.Y(n_216)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_25),
.CON(n_167),
.SN(n_167)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_167),
.A2(n_192),
.B1(n_0),
.B2(n_1),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_89),
.B1(n_87),
.B2(n_71),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_172),
.B1(n_195),
.B2(n_105),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_183),
.B1(n_188),
.B2(n_191),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_114),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_6),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_185),
.C(n_153),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_181),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_133),
.B(n_135),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_144),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_150),
.B1(n_154),
.B2(n_142),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_111),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_186),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_148),
.A2(n_104),
.B1(n_105),
.B2(n_120),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_104),
.B1(n_105),
.B2(n_120),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_142),
.B1(n_156),
.B2(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_186),
.B1(n_189),
.B2(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_223),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_137),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_136),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_146),
.B1(n_96),
.B2(n_139),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_212),
.B1(n_182),
.B2(n_175),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_71),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_139),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_9),
.C(n_14),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_170),
.C(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_9),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_7),
.C(n_13),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_219),
.C(n_180),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_164),
.B(n_190),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_7),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_221),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_15),
.C(n_5),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_5),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_171),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_172),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_218),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_186),
.B1(n_168),
.B2(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_224),
.B1(n_209),
.B2(n_182),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_180),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_175),
.Y(n_263)
);

NOR4xp25_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_223),
.C(n_221),
.D(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_243),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_196),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_210),
.C(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_238),
.C(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_264),
.C(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_251),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_201),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_199),
.B(n_214),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_184),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_184),
.B(n_171),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_5),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_266),
.C(n_229),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_10),
.C(n_11),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_227),
.Y(n_265)
);

XOR2x1_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_12),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_234),
.B1(n_226),
.B2(n_230),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_0),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_246),
.B1(n_239),
.B2(n_231),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_252),
.C(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_253),
.C(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_246),
.B1(n_232),
.B2(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_233),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_287),
.C(n_290),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_266),
.C(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_263),
.C(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_262),
.B1(n_12),
.B2(n_3),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_275),
.B1(n_273),
.B2(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_1),
.C(n_3),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_3),
.B(n_4),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_280),
.B(n_281),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_3),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_294),
.A3(n_284),
.B1(n_287),
.B2(n_290),
.C1(n_283),
.C2(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_271),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_268),
.B(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_302),
.B(n_4),
.Y(n_306)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_4),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_296),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_305),
.Y(n_315)
);

XOR2x1_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_300),
.Y(n_314)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_300),
.B(n_306),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_315),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_312),
.C(n_316),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule