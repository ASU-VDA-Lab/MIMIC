module real_aes_14134_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_781;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_236;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_649;
wire n_162;
wire n_358;
wire n_293;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g325 ( .A(n_0), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_1), .Y(n_165) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_2), .A2(n_49), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g238 ( .A(n_2), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_3), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_4), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_5), .B(n_610), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_6), .B(n_221), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_7), .A2(n_93), .B1(n_136), .B2(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_7), .Y(n_137) );
AND2x2_ASAP7_75t_L g304 ( .A(n_8), .B(n_180), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_9), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_10), .B(n_192), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_11), .B(n_192), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_12), .B(n_611), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_13), .B(n_195), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_14), .B(n_173), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_15), .B(n_324), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_16), .Y(n_687) );
BUFx3_ASAP7_75t_L g157 ( .A(n_17), .Y(n_157) );
INVx1_ASAP7_75t_L g171 ( .A(n_17), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_18), .B(n_179), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_19), .B(n_287), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_20), .Y(n_699) );
BUFx10_ASAP7_75t_L g557 ( .A(n_21), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_22), .B(n_204), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_23), .Y(n_681) );
OAI22x1_ASAP7_75t_SL g575 ( .A1(n_24), .A2(n_78), .B1(n_576), .B2(n_577), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_24), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_25), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_26), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_27), .B(n_610), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_28), .B(n_155), .C(n_339), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_29), .B(n_204), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_30), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_31), .B(n_287), .Y(n_622) );
NAND2xp33_ASAP7_75t_L g640 ( .A(n_32), .B(n_160), .Y(n_640) );
INVx1_ASAP7_75t_L g177 ( .A(n_33), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_34), .A2(n_172), .B(n_289), .C(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_35), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_36), .B(n_167), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_37), .B(n_274), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_38), .B(n_271), .Y(n_654) );
INVx1_ASAP7_75t_L g112 ( .A(n_39), .Y(n_112) );
AND3x2_ASAP7_75t_L g563 ( .A(n_39), .B(n_564), .C(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_40), .B(n_194), .Y(n_193) );
AO221x1_ASAP7_75t_L g607 ( .A1(n_41), .A2(n_83), .B1(n_204), .B2(n_270), .C(n_316), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_42), .B(n_621), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_43), .B(n_169), .Y(n_168) );
AND2x4_ASAP7_75t_L g176 ( .A(n_44), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_45), .B(n_179), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_46), .B(n_188), .Y(n_321) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_47), .B(n_169), .C(n_172), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_48), .B(n_179), .Y(n_212) );
INVx1_ASAP7_75t_L g239 ( .A(n_49), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_50), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_51), .A2(n_295), .B(n_323), .C(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g151 ( .A(n_52), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_53), .A2(n_660), .B(n_662), .C(n_664), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_54), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_55), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g663 ( .A(n_56), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_57), .B(n_188), .Y(n_704) );
AND2x4_ASAP7_75t_L g109 ( .A(n_58), .B(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g255 ( .A(n_59), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_60), .Y(n_911) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_61), .B(n_75), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_62), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_64), .B(n_216), .Y(n_228) );
INVx1_ASAP7_75t_L g269 ( .A(n_65), .Y(n_269) );
AND2x2_ASAP7_75t_L g656 ( .A(n_66), .B(n_188), .Y(n_656) );
INVx1_ASAP7_75t_L g614 ( .A(n_67), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_69), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g128 ( .A(n_69), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_70), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_71), .B(n_159), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_72), .B(n_155), .Y(n_154) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_73), .A2(n_76), .B1(n_610), .B2(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_74), .B(n_172), .Y(n_624) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_77), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g577 ( .A(n_78), .Y(n_577) );
INVx1_ASAP7_75t_L g317 ( .A(n_79), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_80), .B(n_276), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_81), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_82), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g670 ( .A(n_84), .B(n_180), .Y(n_670) );
INVx1_ASAP7_75t_L g163 ( .A(n_85), .Y(n_163) );
BUFx3_ASAP7_75t_L g173 ( .A(n_85), .Y(n_173) );
INVx1_ASAP7_75t_L g198 ( .A(n_85), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_86), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g253 ( .A(n_87), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_88), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_89), .B(n_299), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_90), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_91), .B(n_180), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_92), .B(n_621), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_93), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_94), .B(n_188), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_95), .B(n_226), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_96), .Y(n_248) );
INVx1_ASAP7_75t_L g244 ( .A(n_97), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_98), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_99), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_100), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_117), .B(n_910), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx4f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_104), .Y(n_913) );
OR3x4_ASAP7_75t_SL g104 ( .A(n_105), .B(n_113), .C(n_115), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g580 ( .A(n_111), .Y(n_580) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_112), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_566), .Y(n_117) );
AO21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_554), .B(n_558), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_131), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_120), .A2(n_567), .B(n_573), .Y(n_566) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp67_ASAP7_75t_SL g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_L g564 ( .A(n_128), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_130), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
XNOR2x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_138), .Y(n_134) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_138), .A2(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_480), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_415), .C(n_441), .Y(n_139) );
NAND4xp25_ASAP7_75t_SL g140 ( .A(n_141), .B(n_278), .C(n_371), .D(n_395), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_182), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g543 ( .A(n_143), .Y(n_543) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_144), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g280 ( .A(n_145), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g448 ( .A(n_145), .B(n_357), .Y(n_448) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g354 ( .A(n_146), .B(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g363 ( .A(n_146), .Y(n_363) );
AND2x2_ASAP7_75t_L g472 ( .A(n_146), .B(n_361), .Y(n_472) );
INVx2_ASAP7_75t_L g519 ( .A(n_146), .Y(n_519) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_178), .Y(n_147) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_148), .A2(n_262), .B(n_277), .Y(n_261) );
OAI21x1_ASAP7_75t_L g696 ( .A1(n_148), .A2(n_697), .B(n_704), .Y(n_696) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVxp67_ASAP7_75t_L g631 ( .A(n_149), .Y(n_631) );
BUFx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g240 ( .A(n_151), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_164), .B(n_174), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_158), .B(n_161), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g271 ( .A(n_156), .Y(n_271) );
INVx2_ASAP7_75t_L g610 ( .A(n_156), .Y(n_610) );
INVx2_ASAP7_75t_L g621 ( .A(n_156), .Y(n_621) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_157), .Y(n_218) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
INVx2_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
INVx2_ASAP7_75t_L g265 ( .A(n_160), .Y(n_265) );
INVx3_ASAP7_75t_L g287 ( .A(n_160), .Y(n_287) );
INVx3_ASAP7_75t_L g316 ( .A(n_160), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_161), .A2(n_200), .B(n_202), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_161), .A2(n_273), .B(n_275), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_161), .A2(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g669 ( .A(n_161), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_161), .A2(n_702), .B(n_703), .Y(n_701) );
BUFx10_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g339 ( .A(n_162), .Y(n_339) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g291 ( .A(n_163), .Y(n_291) );
O2A1O1Ixp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_168), .C(n_172), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_166), .A2(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
INVx1_ASAP7_75t_L g227 ( .A(n_170), .Y(n_227) );
INVx2_ASAP7_75t_L g274 ( .A(n_170), .Y(n_274) );
INVx1_ASAP7_75t_L g661 ( .A(n_170), .Y(n_661) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_173), .B(n_246), .Y(n_245) );
NOR3xp33_ASAP7_75t_L g252 ( .A(n_173), .B(n_246), .C(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g270 ( .A(n_173), .Y(n_270) );
INVx1_ASAP7_75t_L g604 ( .A(n_173), .Y(n_604) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_174), .A2(n_333), .B(n_337), .Y(n_332) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_SL g232 ( .A(n_175), .Y(n_232) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_SL g205 ( .A(n_176), .Y(n_205) );
INVx3_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx1_ASAP7_75t_L g303 ( .A(n_176), .Y(n_303) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_179), .Y(n_331) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_207), .Y(n_182) );
OR2x2_ASAP7_75t_L g488 ( .A(n_183), .B(n_311), .Y(n_488) );
AND2x2_ASAP7_75t_L g500 ( .A(n_183), .B(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g385 ( .A(n_184), .Y(n_385) );
AND2x2_ASAP7_75t_L g439 ( .A(n_184), .B(n_368), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_184), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g542 ( .A(n_184), .B(n_424), .Y(n_542) );
AND2x2_ASAP7_75t_L g549 ( .A(n_184), .B(n_209), .Y(n_549) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_185), .Y(n_536) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_206), .Y(n_185) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_186), .A2(n_284), .B(n_362), .Y(n_361) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_186), .A2(n_189), .B(n_206), .Y(n_367) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2x1_ASAP7_75t_SL g230 ( .A(n_187), .B(n_231), .Y(n_230) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g377 ( .A(n_188), .Y(n_377) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_188), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_188), .B(n_246), .Y(n_605) );
INVx2_ASAP7_75t_L g628 ( .A(n_188), .Y(n_628) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_199), .B(n_205), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_197), .Y(n_190) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g201 ( .A(n_195), .Y(n_201) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_195), .Y(n_319) );
INVx2_ASAP7_75t_L g336 ( .A(n_195), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_195), .B(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_196), .Y(n_204) );
INVx2_ASAP7_75t_L g229 ( .A(n_197), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_197), .A2(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g664 ( .A(n_197), .Y(n_664) );
BUFx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx2_ASAP7_75t_L g289 ( .A(n_201), .Y(n_289) );
INVxp67_ASAP7_75t_L g340 ( .A(n_203), .Y(n_340) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_204), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g256 ( .A(n_204), .Y(n_256) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_205), .A2(n_263), .B(n_272), .Y(n_262) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_205), .A2(n_698), .B(n_701), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_207), .A2(n_428), .B(n_483), .C(n_484), .Y(n_482) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_233), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_208), .B(n_453), .Y(n_464) );
OR2x2_ASAP7_75t_L g479 ( .A(n_208), .B(n_456), .Y(n_479) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_208), .Y(n_491) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx2_ASAP7_75t_L g427 ( .A(n_209), .Y(n_427) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g310 ( .A(n_210), .Y(n_310) );
BUFx2_ASAP7_75t_L g345 ( .A(n_210), .Y(n_345) );
OR2x2_ASAP7_75t_L g369 ( .A(n_210), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g374 ( .A(n_210), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g474 ( .A(n_210), .B(n_394), .Y(n_474) );
INVx1_ASAP7_75t_L g531 ( .A(n_210), .Y(n_531) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2x1_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
OAI21x1_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_224), .B(n_230), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_219), .B(n_222), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_216), .A2(n_252), .B1(n_254), .B2(n_256), .Y(n_251) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_217), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g276 ( .A(n_218), .Y(n_276) );
INVx2_ASAP7_75t_L g324 ( .A(n_218), .Y(n_324) );
INVx2_ASAP7_75t_L g611 ( .A(n_218), .Y(n_611) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g297 ( .A(n_222), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_222), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_223), .A2(n_636), .B(n_637), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_228), .B(n_229), .Y(n_224) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_232), .B(n_300), .Y(n_677) );
AND2x2_ASAP7_75t_L g346 ( .A(n_233), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g440 ( .A(n_233), .B(n_433), .Y(n_440) );
AND2x2_ASAP7_75t_L g471 ( .A(n_233), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g505 ( .A(n_233), .Y(n_505) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_259), .Y(n_233) );
INVx1_ASAP7_75t_L g355 ( .A(n_234), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_234), .B(n_517), .Y(n_516) );
AO21x1_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_241), .B(n_257), .Y(n_234) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_235), .A2(n_241), .B(n_257), .Y(n_359) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_236), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_236), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_R g612 ( .A(n_237), .B(n_246), .Y(n_612) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_237) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B1(n_247), .B2(n_249), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_246), .B(n_250), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_246), .B(n_250), .C(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g627 ( .A(n_246), .Y(n_627) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g307 ( .A(n_260), .Y(n_307) );
AND2x2_ASAP7_75t_L g382 ( .A(n_260), .B(n_359), .Y(n_382) );
INVx1_ASAP7_75t_L g391 ( .A(n_260), .Y(n_391) );
INVx1_ASAP7_75t_L g397 ( .A(n_260), .Y(n_397) );
AND2x2_ASAP7_75t_L g409 ( .A(n_260), .B(n_358), .Y(n_409) );
AND2x2_ASAP7_75t_L g444 ( .A(n_260), .B(n_361), .Y(n_444) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_260), .Y(n_463) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B(n_267), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g600 ( .A(n_270), .Y(n_600) );
INVx2_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_308), .B1(n_343), .B2(n_346), .C(n_350), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_305), .Y(n_279) );
AND2x2_ASAP7_75t_L g396 ( .A(n_280), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g413 ( .A(n_282), .B(n_363), .Y(n_413) );
OR2x2_ASAP7_75t_L g430 ( .A(n_282), .B(n_307), .Y(n_430) );
AO31x2_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_298), .A3(n_301), .B(n_304), .Y(n_282) );
AO31x2_ASAP7_75t_L g349 ( .A1(n_283), .A2(n_298), .A3(n_301), .B(n_304), .Y(n_349) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22x1_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_291), .B1(n_292), .B2(n_297), .Y(n_284) );
OAI22x1_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_289), .B2(n_290), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
AOI21x1_ASAP7_75t_L g333 ( .A1(n_291), .A2(n_334), .B(n_335), .Y(n_333) );
AOI21xp5_ASAP7_75t_SL g648 ( .A1(n_291), .A2(n_649), .B(n_650), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_295), .B2(n_296), .Y(n_292) );
AOI21x1_ASAP7_75t_SL g314 ( .A1(n_297), .A2(n_315), .B(n_318), .Y(n_314) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_299), .A2(n_303), .B(n_321), .Y(n_327) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g362 ( .A(n_304), .Y(n_362) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g478 ( .A(n_306), .B(n_460), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_306), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_309), .A2(n_408), .B1(n_410), .B2(n_414), .Y(n_407) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_310), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g399 ( .A(n_310), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_310), .B(n_403), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_310), .B(n_436), .Y(n_435) );
NOR2xp67_ASAP7_75t_R g502 ( .A(n_310), .B(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g384 ( .A(n_311), .B(n_385), .Y(n_384) );
OR2x6_ASAP7_75t_L g311 ( .A(n_312), .B(n_328), .Y(n_311) );
INVx2_ASAP7_75t_L g424 ( .A(n_312), .Y(n_424) );
OR2x2_ASAP7_75t_SL g454 ( .A(n_312), .B(n_375), .Y(n_454) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B(n_327), .Y(n_313) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g402 ( .A(n_328), .B(n_367), .Y(n_402) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_329), .Y(n_370) );
INVx2_ASAP7_75t_L g394 ( .A(n_329), .Y(n_394) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B(n_342), .Y(n_330) );
OA21x2_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_342), .B(n_376), .Y(n_375) );
O2A1O1Ixp5_ASAP7_75t_L g698 ( .A1(n_336), .A2(n_604), .B(n_699), .C(n_700), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_341), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_343), .A2(n_533), .B(n_537), .Y(n_532) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g477 ( .A(n_345), .B(n_439), .Y(n_477) );
OR2x2_ASAP7_75t_L g507 ( .A(n_345), .B(n_393), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_345), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g379 ( .A(n_348), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g389 ( .A(n_348), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g483 ( .A(n_348), .Y(n_483) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g353 ( .A(n_349), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_356), .B(n_364), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_351), .A2(n_387), .B1(n_389), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g381 ( .A(n_353), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_353), .B(n_409), .Y(n_408) );
OR2x6_ASAP7_75t_L g418 ( .A(n_353), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g433 ( .A(n_353), .Y(n_433) );
INVx1_ASAP7_75t_L g419 ( .A(n_354), .Y(n_419) );
INVx1_ASAP7_75t_L g460 ( .A(n_354), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g494 ( .A(n_357), .Y(n_494) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_358), .B(n_363), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_358), .B(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g469 ( .A(n_358), .Y(n_469) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_360), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g468 ( .A(n_360), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g506 ( .A(n_360), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_360), .B(n_382), .Y(n_508) );
AND2x2_ASAP7_75t_L g545 ( .A(n_360), .B(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g517 ( .A(n_361), .Y(n_517) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_369), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_366), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g496 ( .A(n_366), .B(n_427), .Y(n_496) );
INVx1_ASAP7_75t_L g512 ( .A(n_366), .Y(n_512) );
AOI322xp5_ASAP7_75t_L g544 ( .A1(n_366), .A2(n_545), .A3(n_547), .B1(n_549), .B2(n_550), .C1(n_552), .C2(n_553), .Y(n_544) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x4_ASAP7_75t_L g423 ( .A(n_367), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g473 ( .A(n_367), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g485 ( .A(n_367), .B(n_454), .Y(n_485) );
AND2x2_ASAP7_75t_L g388 ( .A(n_368), .B(n_375), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_368), .B(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx1_ASAP7_75t_L g437 ( .A(n_368), .Y(n_437) );
INVx2_ASAP7_75t_L g548 ( .A(n_369), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_378), .B1(n_381), .B2(n_383), .C(n_386), .Y(n_371) );
OR2x2_ASAP7_75t_L g534 ( .A(n_373), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g541 ( .A(n_374), .B(n_542), .Y(n_541) );
OA21x2_ASAP7_75t_L g633 ( .A1(n_376), .A2(n_634), .B(n_641), .Y(n_633) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g429 ( .A(n_380), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g445 ( .A(n_380), .Y(n_445) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
AND2x2_ASAP7_75t_L g537 ( .A(n_382), .B(n_472), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_383), .A2(n_420), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g392 ( .A(n_385), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g450 ( .A(n_387), .Y(n_450) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_390), .Y(n_546) );
INVx2_ASAP7_75t_L g400 ( .A(n_393), .Y(n_400) );
INVx1_ASAP7_75t_L g457 ( .A(n_394), .Y(n_457) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_394), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_401), .B2(n_404), .C(n_407), .Y(n_395) );
INVx2_ASAP7_75t_L g412 ( .A(n_397), .Y(n_412) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_399), .B(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_400), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_401), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g436 ( .A(n_402), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g510 ( .A(n_406), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_409), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_409), .B(n_433), .Y(n_551) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_411), .B(n_494), .Y(n_493) );
NOR2x1p5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g420 ( .A(n_412), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_431), .Y(n_415) );
AOI32xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .A3(n_421), .B1(n_425), .B2(n_428), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g552 ( .A(n_418), .Y(n_552) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g527 ( .A(n_424), .Y(n_527) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g449 ( .A(n_430), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_438), .B2(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_439), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_439), .B(n_474), .Y(n_511) );
INVx1_ASAP7_75t_L g528 ( .A(n_440), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_465), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_447), .B2(n_450), .C(n_451), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g459 ( .A(n_444), .Y(n_459) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_458), .B1(n_461), .B2(n_464), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
AND2x2_ASAP7_75t_L g553 ( .A(n_453), .B(n_549), .Y(n_553) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g529 ( .A(n_454), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OR2x2_ASAP7_75t_L g521 ( .A(n_462), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_473), .B(n_475), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_467), .A2(n_476), .B1(n_478), .B2(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g497 ( .A(n_478), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_520), .C(n_538), .Y(n_480) );
NAND3xp33_ASAP7_75t_SL g481 ( .A(n_482), .B(n_486), .C(n_495), .Y(n_481) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI31xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .A3(n_490), .B(n_492), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g540 ( .A(n_494), .Y(n_540) );
AOI211xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_498), .C(n_509), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_504), .B1(n_507), .B2(n_508), .Y(n_498) );
NOR2xp33_ASAP7_75t_SL g499 ( .A(n_500), .B(n_502), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_500), .B(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_509) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_515), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g523 ( .A(n_519), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_524), .B1(n_528), .B2(n_529), .C(n_532), .Y(n_520) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B(n_544), .Y(n_538) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
CKINVDCx11_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g572 ( .A(n_557), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g571 ( .A(n_564), .B(n_565), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_568), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
BUFx8_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
BUFx8_ASAP7_75t_L g582 ( .A(n_579), .Y(n_582) );
BUFx6f_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_840), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_747), .C(n_783), .D(n_808), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_714), .C(n_730), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_642), .B1(n_689), .B2(n_694), .C(n_705), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_615), .Y(n_589) );
INVx2_ASAP7_75t_L g799 ( .A(n_590), .Y(n_799) );
AND2x4_ASAP7_75t_L g831 ( .A(n_590), .B(n_753), .Y(n_831) );
AND2x2_ASAP7_75t_L g909 ( .A(n_590), .B(n_775), .Y(n_909) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_606), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_591), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g773 ( .A(n_591), .Y(n_773) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_592), .B(n_633), .Y(n_707) );
AND2x2_ASAP7_75t_L g733 ( .A(n_592), .B(n_691), .Y(n_733) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_592), .Y(n_751) );
OR2x2_ASAP7_75t_L g755 ( .A(n_592), .B(n_606), .Y(n_755) );
AND2x2_ASAP7_75t_L g768 ( .A(n_592), .B(n_633), .Y(n_768) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B(n_605), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_600), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_600), .A2(n_684), .B(n_686), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_604), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_604), .A2(n_620), .B(n_622), .Y(n_619) );
OR2x2_ASAP7_75t_L g690 ( .A(n_606), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g708 ( .A(n_606), .B(n_693), .Y(n_708) );
BUFx3_ASAP7_75t_L g721 ( .A(n_606), .Y(n_721) );
INVx2_ASAP7_75t_SL g741 ( .A(n_606), .Y(n_741) );
AND2x2_ASAP7_75t_L g782 ( .A(n_606), .B(n_773), .Y(n_782) );
AND2x2_ASAP7_75t_L g805 ( .A(n_606), .B(n_717), .Y(n_805) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .A3(n_612), .B(n_613), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_611), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g750 ( .A(n_615), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_615), .B(n_772), .Y(n_812) );
AND2x2_ASAP7_75t_L g866 ( .A(n_615), .B(n_741), .Y(n_866) );
AND2x2_ASAP7_75t_L g880 ( .A(n_615), .B(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g846 ( .A(n_616), .B(n_755), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_632), .Y(n_616) );
INVx2_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
BUFx2_ASAP7_75t_SL g729 ( .A(n_617), .Y(n_729) );
AND2x2_ASAP7_75t_L g753 ( .A(n_617), .B(n_633), .Y(n_753) );
INVx1_ASAP7_75t_L g775 ( .A(n_617), .Y(n_775) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
O2A1O1Ixp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_623), .B(n_626), .C(n_629), .Y(n_618) );
INVx2_ASAP7_75t_SL g651 ( .A(n_621), .Y(n_651) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_626), .B(n_648), .Y(n_647) );
AOI21x1_ASAP7_75t_L g652 ( .A1(n_626), .A2(n_653), .B(n_656), .Y(n_652) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_627), .A2(n_635), .B(n_638), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_627), .A2(n_631), .B(n_670), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g691 ( .A(n_633), .Y(n_691) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_633), .Y(n_718) );
INVx1_ASAP7_75t_L g740 ( .A(n_633), .Y(n_740) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_672), .Y(n_642) );
OR2x2_ASAP7_75t_L g722 ( .A(n_643), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g878 ( .A(n_643), .Y(n_878) );
OR2x2_ASAP7_75t_L g902 ( .A(n_643), .B(n_763), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_657), .Y(n_643) );
AND2x2_ASAP7_75t_L g713 ( .A(n_644), .B(n_658), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_644), .B(n_673), .Y(n_795) );
OR2x2_ASAP7_75t_L g824 ( .A(n_644), .B(n_737), .Y(n_824) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g746 ( .A(n_645), .B(n_658), .Y(n_746) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g695 ( .A(n_646), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g727 ( .A(n_646), .Y(n_727) );
AND2x2_ASAP7_75t_L g807 ( .A(n_646), .B(n_738), .Y(n_807) );
OR2x2_ASAP7_75t_L g860 ( .A(n_646), .B(n_658), .Y(n_860) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_647), .B(n_652), .Y(n_646) );
AND2x2_ASAP7_75t_L g736 ( .A(n_657), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g761 ( .A(n_658), .Y(n_761) );
INVx2_ASAP7_75t_L g787 ( .A(n_658), .Y(n_787) );
AND2x2_ASAP7_75t_L g814 ( .A(n_658), .B(n_674), .Y(n_814) );
AO21x2_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_665), .B(n_671), .Y(n_658) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_660), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_661), .B(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B(n_670), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
BUFx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g723 ( .A(n_673), .Y(n_723) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g778 ( .A(n_674), .B(n_779), .Y(n_778) );
OR2x2_ASAP7_75t_L g823 ( .A(n_674), .B(n_787), .Y(n_823) );
INVx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_675), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g829 ( .A(n_675), .B(n_737), .Y(n_829) );
AO21x2_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_682), .Y(n_675) );
AO21x1_ASAP7_75t_SL g712 ( .A1(n_676), .A2(n_678), .B(n_682), .Y(n_712) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
OAI21x1_ASAP7_75t_SL g682 ( .A1(n_677), .A2(n_683), .B(n_688), .Y(n_682) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
OR2x2_ASAP7_75t_L g728 ( .A(n_690), .B(n_729), .Y(n_728) );
NOR2x1_ASAP7_75t_SL g849 ( .A(n_690), .B(n_729), .Y(n_849) );
INVx2_ASAP7_75t_L g792 ( .A(n_692), .Y(n_792) );
INVx2_ASAP7_75t_L g717 ( .A(n_693), .Y(n_717) );
INVx6_ASAP7_75t_L g766 ( .A(n_694), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_694), .B(n_906), .Y(n_905) );
INVx4_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g813 ( .A(n_695), .B(n_814), .Y(n_813) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_695), .Y(n_882) );
INVx2_ASAP7_75t_L g738 ( .A(n_696), .Y(n_738) );
INVxp33_ASAP7_75t_L g779 ( .A(n_696), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVxp67_ASAP7_75t_L g825 ( .A(n_707), .Y(n_825) );
AND2x4_ASAP7_75t_L g732 ( .A(n_708), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g770 ( .A(n_709), .Y(n_770) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .Y(n_709) );
NAND2x1_ASAP7_75t_L g765 ( .A(n_710), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g851 ( .A(n_710), .Y(n_851) );
AND2x2_ASAP7_75t_L g858 ( .A(n_710), .B(n_859), .Y(n_858) );
AND2x4_ASAP7_75t_L g894 ( .A(n_710), .B(n_895), .Y(n_894) );
INVx5_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g785 ( .A(n_711), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g839 ( .A(n_711), .B(n_746), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_711), .B(n_844), .Y(n_843) );
AND2x2_ASAP7_75t_L g865 ( .A(n_711), .B(n_859), .Y(n_865) );
AND2x4_ASAP7_75t_SL g871 ( .A(n_711), .B(n_872), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_711), .B(n_899), .Y(n_898) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g725 ( .A(n_712), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_722), .B1(n_724), .B2(n_728), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
OR2x2_ASAP7_75t_L g833 ( .A(n_716), .B(n_834), .Y(n_833) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g837 ( .A(n_717), .Y(n_837) );
AND2x2_ASAP7_75t_L g900 ( .A(n_717), .B(n_767), .Y(n_900) );
AND2x2_ASAP7_75t_L g818 ( .A(n_718), .B(n_819), .Y(n_818) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g816 ( .A(n_720), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g776 ( .A(n_721), .Y(n_776) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_721), .Y(n_789) );
INVx1_ASAP7_75t_L g834 ( .A(n_721), .Y(n_834) );
AND2x4_ASAP7_75t_L g830 ( .A(n_723), .B(n_746), .Y(n_830) );
OR2x2_ASAP7_75t_L g855 ( .A(n_723), .B(n_806), .Y(n_855) );
OR2x2_ASAP7_75t_L g734 ( .A(n_724), .B(n_735), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND2x4_ASAP7_75t_L g821 ( .A(n_726), .B(n_736), .Y(n_821) );
INVx1_ASAP7_75t_L g845 ( .A(n_726), .Y(n_845) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g899 ( .A(n_727), .B(n_745), .Y(n_899) );
AND2x2_ASAP7_75t_L g885 ( .A(n_729), .B(n_768), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_734), .B1(n_739), .B2(n_742), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_732), .A2(n_871), .B(n_876), .Y(n_875) );
AND2x4_ASAP7_75t_L g804 ( .A(n_733), .B(n_805), .Y(n_804) );
NAND2x1_ASAP7_75t_L g904 ( .A(n_733), .B(n_837), .Y(n_904) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g786 ( .A(n_737), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g745 ( .A(n_738), .Y(n_745) );
INVx1_ASAP7_75t_L g763 ( .A(n_738), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g791 ( .A(n_740), .Y(n_791) );
AOI211x1_ASAP7_75t_L g867 ( .A1(n_740), .A2(n_868), .B(n_873), .C(n_879), .Y(n_867) );
AND2x4_ASAP7_75t_SL g767 ( .A(n_741), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g881 ( .A(n_741), .B(n_773), .Y(n_881) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
AO22x1_ASAP7_75t_L g907 ( .A1(n_743), .A2(n_830), .B1(n_908), .B2(n_909), .Y(n_907) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
OR2x2_ASAP7_75t_L g852 ( .A(n_744), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g870 ( .A(n_744), .Y(n_870) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g874 ( .A(n_745), .B(n_860), .Y(n_874) );
INVx1_ASAP7_75t_L g853 ( .A(n_746), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_756), .B1(n_764), .B2(n_767), .C(n_769), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_752), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI221xp5_ASAP7_75t_SL g783 ( .A1(n_750), .A2(n_784), .B1(n_788), .B2(n_793), .C(n_798), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR2x1_ASAP7_75t_L g862 ( .A(n_755), .B(n_775), .Y(n_862) );
INVx2_ASAP7_75t_L g872 ( .A(n_755), .Y(n_872) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_762), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_760), .Y(n_802) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_SL g895 ( .A(n_763), .B(n_889), .Y(n_895) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g856 ( .A(n_767), .Y(n_856) );
AND2x2_ASAP7_75t_L g810 ( .A(n_768), .B(n_775), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_777), .B2(n_780), .Y(n_769) );
OR2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g848 ( .A(n_772), .Y(n_848) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g819 ( .A(n_773), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g781 ( .A(n_775), .Y(n_781) );
AND2x2_ASAP7_75t_L g908 ( .A(n_775), .B(n_872), .Y(n_908) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g884 ( .A(n_778), .B(n_859), .Y(n_884) );
AND2x2_ASAP7_75t_L g797 ( .A(n_779), .B(n_787), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
INVx1_ASAP7_75t_L g876 ( .A(n_781), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_781), .B(n_782), .Y(n_893) );
AND2x2_ASAP7_75t_L g836 ( .A(n_782), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR2x1_ASAP7_75t_L g864 ( .A(n_786), .B(n_795), .Y(n_864) );
NAND2xp33_ASAP7_75t_L g887 ( .A(n_786), .B(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g828 ( .A(n_787), .Y(n_828) );
AND2x4_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
AND2x4_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_794), .B(n_796), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_796), .A2(n_843), .B(n_846), .C(n_847), .Y(n_842) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B(n_803), .C(n_806), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_815), .C(n_832), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g903 ( .A(n_810), .Y(n_903) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g883 ( .A(n_814), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_820), .B1(n_822), .B2(n_825), .C(n_826), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g906 ( .A(n_823), .Y(n_906) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_830), .B(n_831), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_835), .B(n_838), .Y(n_832) );
INVx1_ASAP7_75t_L g892 ( .A(n_834), .Y(n_892) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
NAND4xp75_ASAP7_75t_L g840 ( .A(n_841), .B(n_867), .C(n_886), .D(n_896), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_850), .B(n_854), .Y(n_841) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_846), .B(n_851), .C(n_852), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_847), .A2(n_874), .B1(n_875), .B2(n_877), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
OAI221xp5_ASAP7_75t_SL g854 ( .A1(n_855), .A2(n_856), .B1(n_857), .B2(n_861), .C(n_863), .Y(n_854) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g889 ( .A(n_860), .Y(n_889) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_862), .A2(n_864), .B1(n_865), .B2(n_866), .Y(n_863) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AO32x1_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_882), .A3(n_883), .B1(n_884), .B2(n_885), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_885), .B(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_890), .B1(n_893), .B2(n_894), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AOI211xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_900), .B(n_901), .C(n_907), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
OAI22xp33_ASAP7_75t_SL g901 ( .A1(n_902), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
endmodule