module real_jpeg_13128_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx1_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_0),
.A2(n_34),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_0),
.B(n_36),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_0),
.A2(n_67),
.B1(n_68),
.B2(n_189),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_0),
.A2(n_68),
.B(n_71),
.C(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_0),
.B(n_93),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_60),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_0),
.B(n_75),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_0),
.A2(n_32),
.B(n_87),
.C(n_296),
.Y(n_295)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_41),
.B1(n_67),
.B2(n_68),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_29),
.B1(n_32),
.B2(n_41),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_41),
.B1(n_56),
.B2(n_62),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_56),
.B1(n_62),
.B2(n_66),
.Y(n_161)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_29),
.B1(n_32),
.B2(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_197),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_7),
.A2(n_56),
.B1(n_62),
.B2(n_197),
.Y(n_281)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_8),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_9),
.A2(n_29),
.B1(n_32),
.B2(n_80),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_80),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_9),
.A2(n_56),
.B1(n_62),
.B2(n_80),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_10),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_134),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_134),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_10),
.A2(n_56),
.B1(n_62),
.B2(n_134),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_12),
.A2(n_29),
.B1(n_32),
.B2(n_170),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_12),
.A2(n_67),
.B1(n_68),
.B2(n_170),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_12),
.A2(n_56),
.B1(n_62),
.B2(n_170),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_38),
.B1(n_56),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_38),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_29),
.B1(n_32),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_86),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_15),
.A2(n_67),
.B1(n_68),
.B2(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_15),
.A2(n_56),
.B1(n_62),
.B2(n_86),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_18),
.A2(n_34),
.B1(n_35),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_18),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_18),
.A2(n_29),
.B1(n_32),
.B2(n_78),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_18),
.A2(n_67),
.B1(n_68),
.B2(n_78),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_18),
.A2(n_56),
.B1(n_62),
.B2(n_78),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_338),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_19),
.B(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B(n_37),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_26),
.A2(n_36),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_26),
.A2(n_36),
.B1(n_40),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_27),
.A2(n_28),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_27),
.A2(n_28),
.B1(n_79),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_28),
.B1(n_77),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_27),
.A2(n_28),
.B1(n_99),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_27),
.A2(n_28),
.B1(n_133),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_27),
.A2(n_28),
.B1(n_196),
.B2(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_29),
.A2(n_32),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_29),
.B(n_189),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_30),
.B(n_32),
.Y(n_187)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_32),
.A2(n_67),
.A3(n_89),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_35),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_39),
.B(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_43),
.B(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_333),
.B(n_335),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_321),
.B(n_332),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_148),
.B(n_318),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_135),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_110),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_49),
.B(n_110),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_81),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_50),
.B(n_96),
.C(n_108),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_76),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_51),
.A2(n_52),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_63),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_54),
.B1(n_76),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_61),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_55),
.A2(n_60),
.B1(n_61),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_55),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_55),
.A2(n_60),
.B1(n_161),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_55),
.A2(n_60),
.B1(n_185),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_55),
.A2(n_60),
.B1(n_225),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_55),
.A2(n_60),
.B1(n_248),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_55),
.A2(n_60),
.B1(n_189),
.B2(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_55),
.A2(n_60),
.B1(n_274),
.B2(n_281),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_56),
.B(n_283),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_124),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_59),
.A2(n_159),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_62),
.A2(n_72),
.B(n_189),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_69),
.B1(n_75),
.B2(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_68),
.B1(n_89),
.B2(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_68),
.B(n_90),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_74),
.B1(n_75),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_75),
.B(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_69),
.A2(n_75),
.B1(n_164),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_69),
.A2(n_75),
.B1(n_213),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_69),
.A2(n_75),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_69),
.A2(n_75),
.B1(n_260),
.B2(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_128),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_73),
.A2(n_165),
.B1(n_240),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_96),
.B1(n_108),
.B2(n_109),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_83),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_94),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_91),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_87),
.A2(n_93),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_87),
.A2(n_93),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_87),
.A2(n_93),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_105),
.B1(n_130),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_91),
.A2(n_130),
.B1(n_131),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_91),
.A2(n_130),
.B1(n_192),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_91),
.A2(n_221),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_98),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_103),
.C(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_98),
.B(n_138),
.C(n_141),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_107),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_106),
.B(n_144),
.C(n_146),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_118),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_132),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_120),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_132),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_135),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_136),
.B(n_137),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_147),
.Y(n_328)
);

OAI21x1_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_173),
.B(n_317),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_171),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_150),
.B(n_171),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_155),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_166),
.C(n_168),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_157),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_162),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_201),
.B(n_316),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_199),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_175),
.B(n_199),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.C(n_181),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_180),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_181),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.C(n_194),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_194),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_232),
.B(n_310),
.C(n_315),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_226),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_203),
.B(n_226),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_216),
.C(n_218),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_204),
.A2(n_205),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_210),
.C(n_215),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_309),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_252),
.B(n_308),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_235),
.B(n_249),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_241),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_302),
.B(n_307),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_290),
.B(n_301),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_270),
.B(n_289),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_256),
.B(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_266),
.C(n_268),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_269),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_278),
.B(n_288),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_276),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_284),
.B(n_287),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_297),
.C(n_299),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_331),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_327),
.B1(n_329),
.B2(n_330),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_329),
.C(n_331),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_334),
.Y(n_337)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule