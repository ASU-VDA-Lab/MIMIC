module fake_jpeg_6495_n_14 (n_3, n_2, n_1, n_0, n_4, n_14);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_14;

wire n_13;
wire n_11;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

NOR2xp33_ASAP7_75t_L g5 ( 
.A(n_3),
.B(n_0),
.Y(n_5)
);

AOI22xp5_ASAP7_75t_L g6 ( 
.A1(n_4),
.A2(n_0),
.B1(n_2),
.B2(n_1),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g7 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_7)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_5),
.B(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_10),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g11 ( 
.A1(n_7),
.A2(n_5),
.B(n_6),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_1),
.B(n_2),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_10),
.B(n_13),
.Y(n_14)
);


endmodule