module fake_jpeg_11195_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_58),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_34),
.B1(n_20),
.B2(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_39),
.B1(n_45),
.B2(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_25),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_22),
.B1(n_43),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_98),
.B1(n_100),
.B2(n_56),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_77),
.B(n_95),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_39),
.B1(n_21),
.B2(n_19),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_39),
.B1(n_21),
.B2(n_19),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_104),
.B1(n_105),
.B2(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_103),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_34),
.B1(n_45),
.B2(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_39),
.B1(n_21),
.B2(n_28),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_48),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_36),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_121),
.B(n_137),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_117),
.B1(n_123),
.B2(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_70),
.A3(n_57),
.B1(n_40),
.B2(n_46),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_46),
.B1(n_45),
.B2(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_45),
.B1(n_46),
.B2(n_68),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_52),
.C(n_46),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_131),
.C(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_130),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_52),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_101),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_38),
.B(n_36),
.C(n_31),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_147),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_85),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_146),
.B(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_166),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_109),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_101),
.B(n_38),
.C(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_159),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_107),
.B(n_38),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_118),
.B(n_133),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_23),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_88),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_77),
.B1(n_111),
.B2(n_120),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_157),
.B1(n_162),
.B2(n_66),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_120),
.B1(n_125),
.B2(n_113),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_122),
.B1(n_118),
.B2(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_31),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_145),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_38),
.B(n_36),
.C(n_25),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_27),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_100),
.B1(n_109),
.B2(n_68),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_66),
.B1(n_36),
.B2(n_93),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_79),
.B1(n_97),
.B2(n_92),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_168),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_129),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_25),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_36),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_171),
.A2(n_183),
.B(n_154),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_177),
.C(n_178),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_189),
.B(n_142),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_184),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_132),
.C(n_130),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_93),
.B1(n_28),
.B2(n_106),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_92),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_106),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_146),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_34),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_167),
.B1(n_164),
.B2(n_36),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_144),
.B1(n_161),
.B2(n_148),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_27),
.C(n_20),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_148),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_202),
.B1(n_204),
.B2(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_197),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_214),
.B1(n_183),
.B2(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_149),
.B1(n_142),
.B2(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_150),
.B1(n_148),
.B2(n_155),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_20),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_218),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_152),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_220),
.C(n_188),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_164),
.B1(n_167),
.B2(n_152),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_171),
.B(n_193),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_27),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_238),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_222),
.B1(n_216),
.B2(n_214),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_201),
.A2(n_193),
.B1(n_190),
.B2(n_196),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_234),
.B1(n_240),
.B2(n_241),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_178),
.C(n_184),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_200),
.C(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_174),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_181),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_189),
.B1(n_180),
.B2(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_202),
.B1(n_204),
.B2(n_207),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_242),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_203),
.B(n_192),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_192),
.B(n_176),
.C(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_194),
.B1(n_176),
.B2(n_20),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_220),
.C(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_219),
.C(n_215),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_255),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_215),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_256),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_227),
.B(n_240),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_9),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_9),
.C(n_1),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_229),
.B1(n_224),
.B2(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_225),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_261),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_10),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_239),
.B(n_241),
.C(n_0),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.C(n_248),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_245),
.A2(n_256),
.B(n_248),
.C(n_255),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

OAI322xp33_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_10),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_267),
.C(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_11),
.C(n_2),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_13),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_12),
.CI(n_4),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_13),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_282),
.B1(n_285),
.B2(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_268),
.C(n_265),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_274),
.A3(n_275),
.B1(n_8),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_277),
.B(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_275),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_271),
.B1(n_268),
.B2(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_265),
.B1(n_5),
.B2(n_14),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_288),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_5),
.C(n_15),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_15),
.C(n_16),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_16),
.B(n_0),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_0),
.Y(n_299)
);


endmodule