module fake_jpeg_1519_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_62),
.Y(n_86)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_59),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_70),
.B(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_61),
.B(n_68),
.C(n_69),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_70),
.CON(n_128),
.SN(n_128)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_84),
.B1(n_67),
.B2(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_76),
.B1(n_57),
.B2(n_72),
.Y(n_122)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_85),
.CI(n_56),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_117),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_53),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_84),
.B1(n_56),
.B2(n_72),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_133),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_8),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_72),
.B1(n_56),
.B2(n_77),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_77),
.B1(n_71),
.B2(n_80),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_63),
.B1(n_60),
.B2(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_0),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_3),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_159),
.C(n_16),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_151),
.B1(n_153),
.B2(n_156),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_142),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_27),
.B1(n_50),
.B2(n_49),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_23),
.B1(n_48),
.B2(n_47),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_24),
.B1(n_45),
.B2(n_42),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_19),
.C(n_40),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_9),
.B(n_10),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_9),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_12),
.B(n_14),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_31),
.B1(n_39),
.B2(n_37),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_14),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_166),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_15),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_17),
.B1(n_28),
.B2(n_34),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_36),
.B(n_51),
.Y(n_175)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_149),
.C(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_158),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_R g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_190),
.Y(n_194)
);

NAND4xp25_ASAP7_75t_SL g187 ( 
.A(n_173),
.B(n_146),
.C(n_167),
.D(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_146),
.CI(n_180),
.CON(n_189),
.SN(n_189)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_179),
.C(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_170),
.B1(n_172),
.B2(n_168),
.Y(n_192)
);

OAI31xp33_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_172),
.A3(n_176),
.B(n_182),
.Y(n_195)
);

BUFx12f_ASAP7_75t_SL g193 ( 
.A(n_191),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_195),
.B(n_190),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_196),
.B(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_188),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_197),
.B(n_186),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_185),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_175),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_187),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_207),
.Y(n_208)
);


endmodule