module fake_jpeg_24258_n_322 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_40),
.B(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_29),
.Y(n_66)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_43),
.B1(n_39),
.B2(n_47),
.Y(n_51)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_31),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_26),
.B1(n_32),
.B2(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_64),
.B(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_28),
.B1(n_24),
.B2(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_28),
.B1(n_36),
.B2(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_18),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_36),
.B1(n_30),
.B2(n_35),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_36),
.B1(n_30),
.B2(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_42),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_54),
.B(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_54),
.B(n_34),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_118),
.Y(n_141)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_58),
.B(n_27),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_68),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_130),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_73),
.B1(n_62),
.B2(n_30),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_121),
.B1(n_86),
.B2(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_128),
.Y(n_169)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_84),
.B1(n_70),
.B2(n_52),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_70),
.B(n_73),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_105),
.B(n_118),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_60),
.B1(n_73),
.B2(n_57),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_87),
.A2(n_100),
.B1(n_106),
.B2(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_57),
.B1(n_50),
.B2(n_80),
.Y(n_139)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_71),
.C(n_80),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_114),
.C(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_97),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_71),
.B1(n_50),
.B2(n_63),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_154),
.B1(n_105),
.B2(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_29),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_123),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_87),
.B(n_20),
.CI(n_74),
.CON(n_153),
.SN(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_91),
.A2(n_50),
.B1(n_27),
.B2(n_23),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_161),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_165),
.C(n_173),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_3),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_132),
.B1(n_149),
.B2(n_143),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_166),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_90),
.C(n_93),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_90),
.Y(n_166)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_125),
.B(n_135),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_93),
.C(n_89),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_137),
.B1(n_153),
.B2(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_88),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_89),
.B1(n_111),
.B2(n_96),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_150),
.B1(n_146),
.B2(n_124),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_101),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_101),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_122),
.B(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_189),
.B(n_171),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_192),
.A2(n_195),
.B(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_182),
.B(n_158),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_152),
.C(n_122),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_197),
.C(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_129),
.C(n_130),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_151),
.C(n_132),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_3),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_207),
.B1(n_155),
.B2(n_175),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_134),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_128),
.B1(n_101),
.B2(n_21),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_88),
.C(n_1),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.C(n_215),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_162),
.C(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_172),
.B1(n_170),
.B2(n_169),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_1),
.C(n_2),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_1),
.B(n_2),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_3),
.C(n_4),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.C(n_5),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_221),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_226),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_240),
.B1(n_214),
.B2(n_191),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_160),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_230),
.B(n_237),
.Y(n_246)
);

NAND5xp2_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_168),
.C(n_186),
.D(n_174),
.E(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_192),
.B1(n_195),
.B2(n_217),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_235),
.B(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_190),
.B(n_183),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_242),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_4),
.B(n_5),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_177),
.B(n_7),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_6),
.B(n_7),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_216),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_230),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_231),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_215),
.B1(n_194),
.B2(n_196),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_194),
.C(n_205),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_257),
.C(n_238),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_218),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_198),
.C(n_8),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_229),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_254),
.C(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_266),
.B(n_269),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_239),
.B(n_222),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_268),
.B(n_273),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_226),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_276),
.Y(n_289)
);

AOI211xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_278),
.B(n_250),
.C(n_230),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_232),
.B1(n_233),
.B2(n_244),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_241),
.B(n_237),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_288),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_252),
.C(n_223),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_243),
.B(n_253),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_262),
.B(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_251),
.B(n_228),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_284),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_276),
.B1(n_257),
.B2(n_228),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_297),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_273),
.B(n_265),
.C(n_255),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_294),
.B1(n_288),
.B2(n_264),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_285),
.B1(n_290),
.B2(n_286),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_291),
.B(n_282),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_261),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_240),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_301),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_309),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_295),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_308),
.B(n_9),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_307),
.B(n_295),
.CI(n_300),
.CON(n_310),
.SN(n_310)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_240),
.A3(n_245),
.B1(n_263),
.B2(n_279),
.C(n_13),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_240),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_313),
.A3(n_306),
.B1(n_303),
.B2(n_305),
.C1(n_14),
.C2(n_10),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_314),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_10),
.C(n_11),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_12),
.A3(n_13),
.B1(n_15),
.B2(n_17),
.C1(n_304),
.C2(n_303),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_311),
.C(n_15),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_318),
.B(n_12),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);


endmodule