module fake_jpeg_11603_n_10 (n_3, n_2, n_1, n_0, n_4, n_10);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_10;

wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

NOR2xp33_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_4),
.Y(n_5)
);

INVx13_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_1),
.B(n_0),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

OAI321xp33_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_9),
.A3(n_5),
.B1(n_6),
.B2(n_2),
.C(n_0),
.Y(n_10)
);

BUFx24_ASAP7_75t_SL g9 ( 
.A(n_7),
.Y(n_9)
);


endmodule