module real_jpeg_27243_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_0),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_289)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_134),
.B(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_30),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_3),
.A2(n_30),
.B(n_160),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_117),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_11),
.B(n_58),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_76),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_96),
.B1(n_97),
.B2(n_211),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_114),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_114),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_114),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_25),
.B1(n_52),
.B2(n_53),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_9),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_10),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_112),
.Y(n_203)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_119),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_119),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_338),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_81),
.B(n_336),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_20),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_21),
.A2(n_43),
.B(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_22),
.A2(n_32),
.B(n_80),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_26),
.B(n_27),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_27),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_23),
.B(n_117),
.CON(n_116),
.SN(n_116)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_32),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_27),
.B(n_30),
.Y(n_131)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_29),
.A2(n_30),
.B1(n_66),
.B2(n_67),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_29),
.A2(n_33),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_29),
.A2(n_52),
.A3(n_65),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_48),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_38),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_73),
.C(n_78),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_39),
.A2(n_40),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_62),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_41),
.A2(n_42),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_43),
.A2(n_48),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_43),
.A2(n_48),
.B1(n_125),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_48),
.B(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_49),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_49),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_49),
.A2(n_62),
.B1(n_304),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_60),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_60),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_50),
.A2(n_57),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_50),
.A2(n_168),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_50),
.A2(n_57),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_50),
.A2(n_57),
.B1(n_167),
.B2(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_50),
.A2(n_57),
.B1(n_91),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_50),
.A2(n_107),
.B(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_53),
.B(n_66),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_53),
.A2(n_56),
.B(n_117),
.C(n_188),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_57),
.B(n_117),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_59),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_61),
.B(n_108),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_62),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_63),
.A2(n_75),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_71),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_64),
.A2(n_71),
.B1(n_111),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_64),
.A2(n_71),
.B1(n_144),
.B2(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_64),
.B(n_70),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_64),
.A2(n_71),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_69),
.A2(n_76),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_75),
.A2(n_77),
.B(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_75),
.A2(n_254),
.B(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_78),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_329),
.B(n_335),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_299),
.A3(n_321),
.B1(n_327),
.B2(n_328),
.C(n_340),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_280),
.B(n_298),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_258),
.B(n_279),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_149),
.B(n_234),
.C(n_257),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_136),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_87),
.B(n_136),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_120),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_104),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_89),
.B(n_104),
.C(n_120),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_90),
.B(n_95),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_92),
.B(n_178),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_98),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_96),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_96),
.A2(n_135),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_96),
.A2(n_135),
.B(n_275),
.Y(n_274)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_97),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_97),
.B(n_117),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_255)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_137),
.A2(n_138),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_142),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_233),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_226),
.B(n_232),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_179),
.B(n_225),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_169),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_153),
.B(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.C(n_165),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_154),
.A2(n_155),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_198),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_176),
.C(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_219),
.B(n_224),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_199),
.B(n_218),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_182),
.B(n_189),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_207),
.B(n_217),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_255),
.B2(n_256),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_246),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_249),
.C(n_253),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_260),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_272),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_267),
.C(n_269),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_274),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_276),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_292),
.B(n_295),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_296),
.B2(n_297),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_291),
.C(n_297),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B(n_290),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_301),
.C(n_311),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_301),
.B1(n_302),
.B2(n_326),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_313),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_308),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_310),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_319),
.C(n_320),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_312),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);


endmodule