module real_aes_9889_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_34;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_39;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_8;
wire n_10;
wire n_33;
wire n_36;
NAND3xp33_ASAP7_75t_SL g14 ( .A(n_0), .B(n_15), .C(n_17), .Y(n_14) );
INVx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
OR2x2_ASAP7_75t_L g34 ( .A(n_1), .B(n_35), .Y(n_34) );
BUFx3_ASAP7_75t_L g32 ( .A(n_2), .Y(n_32) );
INVx1_ASAP7_75t_L g35 ( .A(n_3), .Y(n_35) );
INVx1_ASAP7_75t_L g39 ( .A(n_3), .Y(n_39) );
BUFx2_ASAP7_75t_L g23 ( .A(n_4), .Y(n_23) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_6), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_12), .B1(n_25), .B2(n_33), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
INVx2_ASAP7_75t_L g38 ( .A(n_11), .Y(n_38) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_14), .A2(n_24), .B(n_26), .Y(n_13) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_SL g17 ( .A(n_18), .Y(n_17) );
INVx1_ASAP7_75t_SL g18 ( .A(n_19), .Y(n_18) );
INVx5_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
BUFx8_ASAP7_75t_SL g20 ( .A(n_21), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
BUFx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_27), .Y(n_26) );
INVx1_ASAP7_75t_SL g24 ( .A(n_25), .Y(n_24) );
INVxp67_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
OAI21xp33_ASAP7_75t_L g33 ( .A1(n_28), .A2(n_34), .B(n_36), .Y(n_33) );
INVx1_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
BUFx3_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
AND2x4_ASAP7_75t_L g37 ( .A(n_38), .B(n_39), .Y(n_37) );
endmodule