module real_jpeg_32835_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_526, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_526;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_0),
.Y(n_388)
);

NAND2xp67_ASAP7_75t_SL g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_1),
.B(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_1),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_1),
.B(n_510),
.Y(n_509)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.A3(n_482),
.B1(n_521),
.B2(n_523),
.C(n_526),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_2),
.B(n_522),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_6),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_6),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_6),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_6),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_6),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_50),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_7),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_155),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_7),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_8),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_8),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_8),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_9),
.B(n_249),
.Y(n_248)
);

NAND2x1_ASAP7_75t_L g263 ( 
.A(n_9),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_9),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_9),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_9),
.B(n_422),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_10),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_11),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_103),
.Y(n_161)
);

NAND2x2_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_13),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_14),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_14),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_14),
.B(n_54),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_14),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_14),
.B(n_255),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_14),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_14),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_14),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_15),
.Y(n_403)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_17),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_17),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_17),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_17),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_17),
.B(n_399),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_17),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_19),
.B(n_524),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_205),
.B(n_480),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_22),
.B(n_166),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_91),
.C(n_126),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_23),
.B(n_92),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_60),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_24),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.C(n_47),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_25),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_35),
.C(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_31),
.A2(n_95),
.B1(n_104),
.B2(n_105),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_31),
.A2(n_73),
.B1(n_154),
.B2(n_312),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g431 ( 
.A1(n_34),
.A2(n_35),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_44),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_35),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_35),
.B(n_435),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_38),
.B(n_47),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_46),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_42),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_44),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_44),
.A2(n_144),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_44),
.B(n_222),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_45),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_45),
.Y(n_411)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_45),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_46),
.B(n_243),
.C(n_248),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_46),
.B(n_466),
.Y(n_465)
);

XNOR2x1_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_49),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_49),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_49),
.B(n_198),
.C(n_262),
.Y(n_298)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_51),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_56),
.C(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_55),
.Y(n_199)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_74),
.B2(n_90),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_61),
.Y(n_169)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_64),
.A2(n_71),
.B1(n_87),
.B2(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_64),
.B(n_69),
.C(n_72),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_64),
.A2(n_71),
.B1(n_495),
.B2(n_498),
.Y(n_494)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_75),
.C(n_86),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_75),
.B(n_163),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_83),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_76),
.A2(n_83),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_76),
.A2(n_130),
.B1(n_176),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_76),
.B(n_181),
.C(n_182),
.Y(n_500)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_82),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_82),
.Y(n_397)
);

CKINVDCx12_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_89),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_106),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_94),
.B(n_108),
.C(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_96),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_96),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_96),
.B(n_99),
.C(n_104),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_96),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_96),
.B(n_213),
.C(n_215),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_96),
.A2(n_223),
.B(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_96),
.B(n_198),
.Y(n_516)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_98),
.Y(n_297)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_98),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_125),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_133),
.C(n_137),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_113),
.B(n_119),
.C(n_121),
.Y(n_202)
);

HB1xp67_ASAP7_75t_SL g300 ( 
.A(n_113),
.Y(n_300)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_115),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_124),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_124),
.Y(n_275)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_124),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_126),
.B(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_145),
.B(n_165),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_127),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_141),
.Y(n_127)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_128),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_132),
.A2(n_141),
.B1(n_142),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_132),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_133),
.A2(n_137),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_133),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_133),
.A2(n_303),
.B1(n_504),
.B2(n_506),
.Y(n_503)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_135),
.Y(n_422)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_137),
.Y(n_302)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_162),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_162),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_146),
.B(n_162),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_158),
.C(n_161),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_147),
.A2(n_148),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_154),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_149),
.B(n_151),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_154),
.Y(n_312)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_160),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_161),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_167),
.B(n_486),
.C(n_487),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_172),
.B(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_173),
.B(n_174),
.C(n_518),
.Y(n_517)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_187),
.Y(n_518)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_188),
.Y(n_488)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_189),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_190),
.B(n_202),
.C(n_203),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI21x1_ASAP7_75t_SL g513 ( 
.A1(n_192),
.A2(n_514),
.B(n_516),
.Y(n_513)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_197),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_198),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_361),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_339),
.B(n_353),
.C(n_360),
.Y(n_206)
);

AOI21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_314),
.B(n_338),
.Y(n_207)
);

NAND2x1p5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_288),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g363 ( 
.A(n_209),
.B(n_288),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_240),
.C(n_266),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_211),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.C(n_226),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_212),
.B(n_460),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_219),
.A2(n_220),
.B1(n_226),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_225),
.Y(n_378)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_226),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.C(n_235),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_227),
.A2(n_228),
.B1(n_235),
.B2(n_236),
.Y(n_450)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_231),
.B(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_241),
.B(n_267),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_242),
.B(n_253),
.C(n_260),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_243),
.B(n_248),
.Y(n_466)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_257),
.B(n_259),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_257),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_330),
.C(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_283),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_284),
.C(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_276),
.C(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_280),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_305),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_306),
.C(n_307),
.Y(n_337)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_304),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_299),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_304),
.C(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_294),
.C(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_337),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_341),
.C(n_342),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_332),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_319),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_328),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_338),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_343),
.B1(n_354),
.B2(n_358),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_340),
.B(n_343),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_344),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.C(n_347),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_349),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_358),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_354),
.B(n_358),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.C(n_357),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_475),
.C(n_476),
.Y(n_361)
);

NOR2x1p5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_469),
.B(n_474),
.Y(n_364)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_457),
.B(n_468),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_437),
.B(n_455),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_413),
.B(n_436),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_390),
.B(n_412),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_385),
.B(n_389),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_376),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_379),
.B1(n_380),
.B2(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_379),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_384),
.Y(n_391)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_407),
.Y(n_406)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_392),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_404),
.B2(n_405),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_398),
.C(n_404),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_408),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_424),
.Y(n_423)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_415),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_427),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_428),
.C(n_431),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_423),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_421),
.C(n_423),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_432),
.Y(n_435)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_451),
.C(n_454),
.Y(n_437)
);

O2A1O1Ixp5_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_439),
.B(n_454),
.C(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_445),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_439),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_444),
.C(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_448),
.C(n_452),
.Y(n_467)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_453),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_467),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_467),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_463),
.C(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_465),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_465),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_472),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_479),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_521),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_519),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_489),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_489),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_517),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_502),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_493)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_507),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_505),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_512),
.B2(n_513),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);


endmodule