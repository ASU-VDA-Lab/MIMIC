module fake_jpeg_22275_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_20),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_8),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_14),
.B1(n_9),
.B2(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_29),
.B(n_18),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_12),
.B1(n_9),
.B2(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_36),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_11),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_23),
.Y(n_39)
);

AND2x6_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_3),
.Y(n_42)
);

A2O1A1O1Ixp25_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_4),
.B(n_5),
.C(n_13),
.D(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_30),
.B1(n_26),
.B2(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_34),
.CI(n_38),
.CON(n_48),
.SN(n_48)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_49),
.B(n_4),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_49),
.C(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_53),
.B(n_54),
.C(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_54),
.Y(n_58)
);


endmodule