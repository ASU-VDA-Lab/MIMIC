module fake_jpeg_16570_n_92 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_0),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_55),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_45),
.B1(n_36),
.B2(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_41),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_62),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_76),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_68),
.B(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_7),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_80),
.B1(n_11),
.B2(n_14),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_9),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_15),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_17),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_21),
.B(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_27),
.B(n_29),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_30),
.CI(n_31),
.CON(n_92),
.SN(n_92)
);


endmodule