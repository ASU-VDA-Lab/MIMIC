module fake_jpeg_20400_n_295 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_295);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_31),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_21),
.B1(n_17),
.B2(n_25),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_35),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_33),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_65),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_34),
.Y(n_74)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_78),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_32),
.B(n_33),
.C(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_72),
.B1(n_42),
.B2(n_49),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_36),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_74),
.B(n_80),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_36),
.B1(n_42),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_40),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_40),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_34),
.C(n_44),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_70),
.B1(n_83),
.B2(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_20),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_100),
.Y(n_121)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_68),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_34),
.C(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_20),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_18),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_18),
.B(n_24),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_55),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_85),
.B(n_83),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_28),
.B1(n_94),
.B2(n_34),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_71),
.B(n_74),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_112),
.B(n_84),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_28),
.B1(n_81),
.B2(n_25),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_72),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_101),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_74),
.B1(n_78),
.B2(n_80),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_116),
.B1(n_39),
.B2(n_96),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_74),
.B1(n_80),
.B2(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_50),
.B1(n_76),
.B2(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_69),
.B1(n_81),
.B2(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_59),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_149),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_97),
.C(n_87),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_115),
.C(n_123),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_132),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_87),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_67),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_150),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_64),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_146),
.B1(n_130),
.B2(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_126),
.B1(n_105),
.B2(n_81),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_112),
.B(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_107),
.B(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_79),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_144),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_176),
.B(n_113),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_182),
.C(n_183),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_131),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_168),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_147),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_167),
.C(n_169),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_105),
.B(n_112),
.C(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_153),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_132),
.B(n_120),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_60),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_130),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_79),
.C(n_68),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_154),
.C(n_153),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_196),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_190),
.B(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_143),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_168),
.B(n_175),
.C(n_164),
.D(n_163),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_190),
.B(n_184),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_162),
.B1(n_160),
.B2(n_173),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_203),
.B1(n_206),
.B2(n_28),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_51),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_201),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_176),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_55),
.C(n_60),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_184),
.C(n_193),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_21),
.B1(n_39),
.B2(n_17),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_223),
.C(n_206),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_171),
.B1(n_157),
.B2(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_216),
.B1(n_203),
.B2(n_202),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_159),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_224),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_188),
.B1(n_166),
.B2(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_216),
.B1(n_220),
.B2(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_225),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_59),
.B1(n_29),
.B2(n_11),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_195),
.B(n_196),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_55),
.C(n_60),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_192),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_12),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_195),
.B1(n_59),
.B2(n_2),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_234),
.B1(n_238),
.B2(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_15),
.B(n_23),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_10),
.B(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_19),
.B1(n_15),
.B2(n_23),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_241),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_211),
.C(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_217),
.C(n_225),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_248),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_226),
.B1(n_237),
.B2(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.C(n_254),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_217),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_250),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_62),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_228),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_252),
.B(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_262),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.C(n_34),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_234),
.C(n_62),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_62),
.C(n_56),
.Y(n_263)
);

AOI221xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_12),
.B1(n_56),
.B2(n_4),
.C(n_5),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_12),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_258),
.C(n_257),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_275),
.B(n_3),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_9),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_56),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_16),
.C(n_14),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_29),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_14),
.C(n_4),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_14),
.C(n_5),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_3),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_283),
.B(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_277),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_286),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_270),
.B(n_267),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_5),
.B(n_6),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_6),
.C(n_7),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_6),
.B(n_7),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_7),
.B(n_8),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_8),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_8),
.B(n_9),
.Y(n_295)
);


endmodule