module fake_jpeg_26689_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_17),
.B(n_31),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_8),
.C(n_14),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_61),
.B1(n_64),
.B2(n_39),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_44),
.B1(n_42),
.B2(n_19),
.Y(n_87)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_82),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_97),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_30),
.B1(n_17),
.B2(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_73),
.B1(n_83),
.B2(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_39),
.B1(n_36),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_99),
.B1(n_101),
.B2(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_90),
.B(n_93),
.C(n_35),
.Y(n_131)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_16),
.B1(n_35),
.B2(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_85),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_89),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_18),
.B1(n_23),
.B2(n_36),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_25),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_25),
.Y(n_92)
);

OR2x4_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_16),
.Y(n_93)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_16),
.B1(n_21),
.B2(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_24),
.B1(n_21),
.B2(n_35),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_42),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_21),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_19),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_27),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_27),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_130),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_126),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_40),
.B1(n_36),
.B2(n_59),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_117),
.B1(n_76),
.B2(n_77),
.Y(n_147)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_20),
.B1(n_23),
.B2(n_18),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_135),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_89),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_40),
.C(n_36),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_115),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_126),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_91),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_116),
.B1(n_115),
.B2(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_158),
.B1(n_125),
.B2(n_110),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_137),
.B(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_80),
.B(n_85),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_145),
.B(n_159),
.Y(n_179)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_148),
.B1(n_149),
.B2(n_19),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_146),
.Y(n_188)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_163),
.B1(n_164),
.B2(n_68),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_160),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_166),
.B1(n_133),
.B2(n_97),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_127),
.B1(n_96),
.B2(n_34),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_154),
.B(n_7),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_40),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_95),
.B1(n_68),
.B2(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_75),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_75),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_165),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_106),
.B1(n_69),
.B2(n_77),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_113),
.A2(n_122),
.B1(n_110),
.B2(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_105),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_174),
.B1(n_194),
.B2(n_144),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_121),
.C(n_125),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_182),
.C(n_189),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_183),
.B1(n_185),
.B2(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_84),
.B1(n_81),
.B2(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_150),
.B(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_175),
.B(n_176),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_118),
.B1(n_100),
.B2(n_96),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_145),
.B1(n_166),
.B2(n_147),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_154),
.C(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_118),
.B1(n_133),
.B2(n_22),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_42),
.C(n_23),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_138),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_20),
.A3(n_22),
.B1(n_18),
.B2(n_23),
.C1(n_11),
.C2(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_187),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_34),
.B1(n_18),
.B2(n_20),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_137),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_141),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_139),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_186),
.B1(n_190),
.B2(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_210),
.B1(n_219),
.B2(n_178),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_178),
.B(n_184),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_156),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_167),
.B1(n_152),
.B2(n_149),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_146),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_221),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_15),
.C(n_2),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_1),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_10),
.C(n_14),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_195),
.C(n_196),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_179),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_242),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_179),
.C(n_181),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.C(n_235),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_191),
.C(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_243),
.B1(n_206),
.B2(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_6),
.C(n_13),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_6),
.C(n_13),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_239),
.C(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_15),
.C(n_12),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_11),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_207),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_1),
.B(n_2),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_250),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_256),
.B(n_200),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_203),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_259),
.B(n_230),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_219),
.B1(n_216),
.B2(n_198),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_257),
.B1(n_210),
.B2(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_213),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_246),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_223),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_244),
.B1(n_251),
.B2(n_227),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_225),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_271),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_229),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_274),
.C(n_258),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_256),
.B1(n_244),
.B2(n_227),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_209),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_2),
.B(n_3),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_266),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_241),
.B1(n_212),
.B2(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_222),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_224),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_211),
.B1(n_208),
.B2(n_238),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_285),
.B1(n_267),
.B2(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_265),
.B(n_261),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_284),
.C(n_280),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_298),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_276),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_287),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_294),
.C(n_295),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_288),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_299),
.B(n_286),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_274),
.B(n_4),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_5),
.B(n_3),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_3),
.C(n_4),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_4),
.Y(n_308)
);


endmodule