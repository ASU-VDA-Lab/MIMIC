module fake_jpeg_499_n_402 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_402);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_402;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_58),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g169 ( 
.A(n_60),
.Y(n_169)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_7),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_64),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_71),
.Y(n_132)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_68),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_54),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_78),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_76),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_28),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_81),
.B(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_17),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_31),
.B(n_0),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_99),
.B(n_102),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_33),
.B(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_33),
.B(n_15),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_42),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_43),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_111),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_42),
.B(n_16),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_16),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_115),
.B(n_139),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_27),
.B1(n_38),
.B2(n_48),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_125),
.A2(n_128),
.B1(n_147),
.B2(n_173),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_25),
.B1(n_43),
.B2(n_27),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_135),
.B(n_158),
.Y(n_187)
);

OA22x2_ASAP7_75t_SL g137 ( 
.A1(n_83),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_137),
.A2(n_152),
.B1(n_161),
.B2(n_119),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_84),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_48),
.B1(n_0),
.B2(n_17),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_144),
.B1(n_148),
.B2(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_165),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_0),
.B1(n_16),
.B2(n_86),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_80),
.B1(n_85),
.B2(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_146),
.A2(n_159),
.B1(n_170),
.B2(n_172),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_97),
.B1(n_105),
.B2(n_94),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_87),
.A2(n_90),
.B1(n_108),
.B2(n_96),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_91),
.A2(n_73),
.B1(n_66),
.B2(n_107),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_77),
.B1(n_64),
.B2(n_112),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_76),
.C(n_56),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_123),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_68),
.B(n_98),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_76),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_56),
.A2(n_88),
.B(n_71),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_182),
.B(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_93),
.B(n_63),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_89),
.A2(n_18),
.B1(n_38),
.B2(n_37),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_89),
.A2(n_18),
.B1(n_38),
.B2(n_37),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_74),
.A2(n_79),
.B1(n_89),
.B2(n_101),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_63),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_63),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_71),
.A2(n_104),
.B(n_63),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_121),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_214),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_198),
.Y(n_252)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_194),
.B(n_211),
.Y(n_267)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_169),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_196),
.B(n_215),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_128),
.A2(n_173),
.B1(n_149),
.B2(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_197),
.A2(n_241),
.B1(n_240),
.B2(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_199),
.B(n_202),
.Y(n_259)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_123),
.B(n_125),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_142),
.B(n_129),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_205),
.Y(n_269)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_130),
.B(n_134),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_206),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_116),
.B(n_131),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_208),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_123),
.B(n_183),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_214),
.C(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_117),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_218),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_141),
.B(n_177),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_156),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_145),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_137),
.A2(n_181),
.B1(n_162),
.B2(n_154),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_225),
.B1(n_120),
.B2(n_233),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_124),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_223),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_118),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_136),
.B(n_163),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_137),
.A2(n_118),
.B1(n_119),
.B2(n_155),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_230),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_122),
.B(n_127),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_147),
.B(n_155),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_126),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_152),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_237),
.Y(n_280)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_127),
.B(n_171),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_167),
.B1(n_133),
.B2(n_120),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_240),
.B(n_208),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_167),
.A2(n_125),
.B1(n_123),
.B2(n_74),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_133),
.A2(n_160),
.B1(n_146),
.B2(n_79),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_120),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_196),
.B1(n_211),
.B2(n_235),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_265),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_188),
.B(n_224),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_246),
.A2(n_277),
.B(n_256),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_201),
.C(n_194),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_261),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_187),
.B(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_281),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_254),
.A2(n_263),
.B1(n_245),
.B2(n_255),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_268),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_201),
.A2(n_209),
.B1(n_217),
.B2(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_256),
.A2(n_265),
.B1(n_268),
.B2(n_272),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_210),
.A2(n_224),
.B1(n_228),
.B2(n_192),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_228),
.B1(n_186),
.B2(n_220),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_238),
.B1(n_239),
.B2(n_202),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_185),
.A2(n_193),
.B(n_204),
.C(n_229),
.Y(n_270)
);

HAxp5_ASAP7_75t_SL g302 ( 
.A(n_270),
.B(n_269),
.CON(n_302),
.SN(n_302)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_195),
.A2(n_200),
.B1(n_216),
.B2(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_231),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_237),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_191),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_283),
.B(n_286),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_212),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_306),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_288),
.B(n_308),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_249),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_294),
.B(n_300),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_266),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_293),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_277),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_297),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_314),
.B1(n_274),
.B2(n_262),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_304),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_310),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_272),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_245),
.B(n_258),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_248),
.B(n_247),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_250),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_307),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_280),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_261),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_273),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_244),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_261),
.CI(n_251),
.CON(n_315),
.SN(n_315)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_315),
.A2(n_331),
.B(n_300),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_267),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_322),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_267),
.C(n_276),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_326),
.A2(n_294),
.B(n_303),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_247),
.C(n_270),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_332),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_279),
.C(n_275),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_286),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_313),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_275),
.C(n_257),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_333),
.B(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_314),
.B1(n_288),
.B2(n_296),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_332),
.C(n_326),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_333),
.B(n_308),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_295),
.Y(n_349)
);

HAxp5_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_351),
.CON(n_360),
.SN(n_360)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_319),
.B(n_284),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_327),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_353),
.B(n_285),
.Y(n_357)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_312),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_354),
.A2(n_337),
.B1(n_335),
.B2(n_328),
.Y(n_356)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_367),
.C(n_344),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_322),
.C(n_316),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_375),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_299),
.B1(n_289),
.B2(n_317),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_377),
.Y(n_384)
);

OA21x2_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_338),
.B(n_349),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_374),
.B(n_376),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_366),
.B(n_342),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_321),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_298),
.B1(n_352),
.B2(n_299),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_284),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_SL g376 ( 
.A(n_361),
.B(n_340),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_342),
.C(n_346),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_369),
.C(n_373),
.Y(n_380)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_363),
.A3(n_355),
.B1(n_358),
.B2(n_341),
.C1(n_354),
.C2(n_362),
.Y(n_379)
);

AOI21xp33_ASAP7_75t_L g392 ( 
.A1(n_379),
.A2(n_337),
.B(n_320),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_380),
.B(n_383),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_362),
.C(n_336),
.Y(n_383)
);

AOI31xp67_ASAP7_75t_SL g385 ( 
.A1(n_371),
.A2(n_329),
.A3(n_360),
.B(n_323),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_386),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_384),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_392),
.B(n_368),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_357),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g396 ( 
.A1(n_390),
.A2(n_391),
.B(n_318),
.C(n_294),
.Y(n_396)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_377),
.A3(n_317),
.B1(n_370),
.B2(n_368),
.C1(n_289),
.C2(n_356),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_394),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_380),
.C(n_383),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_382),
.B(n_386),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_396),
.C(n_323),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_364),
.B(n_353),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_399),
.A2(n_400),
.B(n_290),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_364),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_345),
.Y(n_402)
);


endmodule