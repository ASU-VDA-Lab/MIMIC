module fake_jpeg_12063_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_282;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_40),
.B(n_61),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_22),
.A2(n_7),
.B(n_1),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_4),
.B(n_9),
.C(n_11),
.Y(n_99)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_58),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_83),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_20),
.B1(n_27),
.B2(n_37),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_32),
.B1(n_20),
.B2(n_27),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_20),
.B1(n_27),
.B2(n_35),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_17),
.B1(n_35),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_19),
.B1(n_17),
.B2(n_35),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_76),
.B1(n_82),
.B2(n_86),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_19),
.B1(n_17),
.B2(n_16),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_37),
.B1(n_36),
.B2(n_26),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_19),
.B1(n_31),
.B2(n_30),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_60),
.B1(n_59),
.B2(n_47),
.Y(n_80)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_21),
.B1(n_16),
.B2(n_0),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_81),
.A2(n_80),
.B(n_94),
.C(n_87),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_33),
.B1(n_25),
.B2(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_26),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_60),
.B1(n_59),
.B2(n_46),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_29),
.B1(n_21),
.B2(n_0),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_43),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_13),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_15),
.B1(n_42),
.B2(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_15),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_68),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_71),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_111),
.B(n_129),
.Y(n_158)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_124),
.Y(n_169)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_137),
.B1(n_122),
.B2(n_107),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_99),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_86),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_106),
.Y(n_136)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_97),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_71),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_97),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_116),
.B1(n_123),
.B2(n_141),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_81),
.B1(n_78),
.B2(n_95),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_153),
.B1(n_161),
.B2(n_157),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_81),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_78),
.B1(n_95),
.B2(n_74),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_130),
.A3(n_119),
.B1(n_127),
.B2(n_112),
.Y(n_154)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_162),
.A3(n_151),
.B(n_153),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_94),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_74),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_155),
.C(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_66),
.B1(n_134),
.B2(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_167),
.B1(n_168),
.B2(n_175),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_66),
.B1(n_108),
.B2(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_128),
.B1(n_109),
.B2(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_127),
.B1(n_113),
.B2(n_120),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_144),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_137),
.B1(n_139),
.B2(n_107),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_131),
.B1(n_115),
.B2(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_162),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_186),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_194),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_144),
.B1(n_152),
.B2(n_202),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_187),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_158),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_143),
.B(n_150),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_198),
.B(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_145),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_202),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_154),
.B(n_148),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_161),
.B(n_156),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_170),
.B(n_167),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_203),
.B(n_204),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_147),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_155),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_228),
.B1(n_206),
.B2(n_199),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_183),
.B(n_200),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_224),
.B(n_227),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_152),
.B(n_208),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_198),
.B(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_180),
.B1(n_203),
.B2(n_193),
.Y(n_228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_204),
.B(n_189),
.C(n_190),
.D(n_181),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_209),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_181),
.A2(n_195),
.B1(n_179),
.B2(n_197),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_179),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_218),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_244),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_213),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_242),
.B1(n_243),
.B2(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_241),
.B(n_246),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_212),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.C(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_227),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_231),
.B(n_233),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_251),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_231),
.B(n_224),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_222),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_220),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_215),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_252),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_211),
.B1(n_216),
.B2(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_260),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_230),
.B1(n_220),
.B2(n_221),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_239),
.B1(n_253),
.B2(n_251),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_249),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_235),
.B1(n_243),
.B2(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_248),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_257),
.C(n_263),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_257),
.B(n_259),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_260),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_271),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_244),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_262),
.CI(n_261),
.CON(n_276),
.SN(n_276)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_262),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_254),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_271),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_285),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_283),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_259),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_286),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.B(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_297),
.A3(n_288),
.B1(n_289),
.B2(n_273),
.C(n_274),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_258),
.B(n_281),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_302),
.Y(n_303)
);


endmodule