module real_aes_6517_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_725, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_725;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_0), .A2(n_180), .B(n_181), .C(n_185), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_1), .B(n_174), .Y(n_187) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_3), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_4), .A2(n_148), .B(n_165), .C(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_168), .B(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_6), .A2(n_168), .B(n_270), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_7), .A2(n_37), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_7), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_7), .B(n_174), .Y(n_500) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_8), .A2(n_140), .B(n_227), .Y(n_226) );
AND2x6_ASAP7_75t_L g165 ( .A(n_9), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_10), .A2(n_148), .B(n_165), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g465 ( .A(n_11), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_12), .B(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_12), .B(n_43), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_13), .B(n_184), .Y(n_475) );
INVx1_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_15), .B(n_159), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_16), .B(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_17), .A2(n_160), .B(n_484), .C(n_486), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_18), .B(n_174), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_19), .A2(n_68), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_19), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_20), .B(n_217), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_21), .A2(n_148), .B(n_211), .C(n_216), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_22), .A2(n_183), .B(n_235), .C(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_23), .B(n_184), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_24), .B(n_184), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_25), .Y(n_503) );
INVx1_ASAP7_75t_L g515 ( .A(n_26), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_27), .A2(n_148), .B(n_216), .C(n_230), .Y(n_229) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_29), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_30), .A2(n_436), .B1(n_705), .B2(n_706), .C1(n_715), .C2(n_718), .Y(n_435) );
INVx1_ASAP7_75t_L g532 ( .A(n_31), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_32), .A2(n_168), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g150 ( .A(n_33), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_34), .A2(n_163), .B(n_195), .C(n_196), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_35), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_36), .A2(n_183), .B(n_497), .C(n_499), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_37), .Y(n_128) );
INVxp67_ASAP7_75t_L g533 ( .A(n_38), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_39), .B(n_232), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_40), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_41), .A2(n_148), .B(n_216), .C(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_42), .A2(n_105), .B1(n_118), .B2(n_723), .Y(n_104) );
INVx1_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_44), .A2(n_185), .B(n_463), .C(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_45), .B(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_46), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_47), .B(n_159), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_48), .B(n_168), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_49), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_50), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_51), .A2(n_163), .B(n_195), .C(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_SL g706 ( .A1(n_52), .A2(n_707), .B1(n_708), .B2(n_714), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_52), .Y(n_714) );
INVx1_ASAP7_75t_L g182 ( .A(n_53), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_54), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_54), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_55), .A2(n_85), .B1(n_712), .B2(n_713), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_55), .Y(n_713) );
INVx1_ASAP7_75t_L g257 ( .A(n_56), .Y(n_257) );
INVx1_ASAP7_75t_L g453 ( .A(n_57), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_58), .B(n_168), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_59), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g461 ( .A(n_60), .Y(n_461) );
INVx1_ASAP7_75t_L g166 ( .A(n_61), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_62), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_63), .B(n_174), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_64), .A2(n_155), .B(n_215), .C(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
INVx1_ASAP7_75t_SL g498 ( .A(n_66), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_67), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_68), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_69), .B(n_159), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_70), .B(n_174), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_71), .B(n_160), .Y(n_246) );
INVx1_ASAP7_75t_L g506 ( .A(n_72), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_73), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_74), .B(n_199), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_75), .A2(n_148), .B(n_153), .C(n_163), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_76), .Y(n_271) );
INVx1_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_78), .A2(n_168), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_79), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_80), .A2(n_168), .B(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_81), .A2(n_209), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g482 ( .A(n_82), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_83), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_84), .B(n_198), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_85), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_86), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_87), .A2(n_168), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g485 ( .A(n_88), .Y(n_485) );
INVx2_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
INVx1_ASAP7_75t_L g474 ( .A(n_90), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_91), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_92), .B(n_184), .Y(n_247) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_93), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g428 ( .A(n_93), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g439 ( .A(n_93), .B(n_430), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_93), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_94), .A2(n_148), .B(n_163), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_95), .B(n_168), .Y(n_193) );
INVx1_ASAP7_75t_L g197 ( .A(n_96), .Y(n_197) );
INVxp67_ASAP7_75t_L g274 ( .A(n_97), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_98), .B(n_140), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g154 ( .A(n_100), .Y(n_154) );
INVx1_ASAP7_75t_L g242 ( .A(n_101), .Y(n_242) );
INVx2_ASAP7_75t_L g456 ( .A(n_102), .Y(n_456) );
AND2x2_ASAP7_75t_L g259 ( .A(n_103), .B(n_202), .Y(n_259) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx5_ASAP7_75t_SL g723 ( .A(n_108), .Y(n_723) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_115), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g430 ( .A(n_111), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AO21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_434), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g722 ( .A(n_121), .Y(n_722) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_426), .B(n_432), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_424), .B2(n_425), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_126), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_129), .Y(n_425) );
XNOR2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_133), .Y(n_129) );
INVx2_ASAP7_75t_L g440 ( .A(n_133), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_133), .A2(n_438), .B1(n_720), .B2(n_721), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_367), .Y(n_133) );
AND4x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_307), .C(n_322), .D(n_347), .Y(n_134) );
NOR2xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_280), .Y(n_135) );
OAI21xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_188), .B(n_260), .Y(n_136) );
AND2x2_ASAP7_75t_L g310 ( .A(n_137), .B(n_206), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_137), .B(n_205), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_137), .B(n_189), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_137), .Y(n_377) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_173), .Y(n_137) );
INVx2_ASAP7_75t_L g294 ( .A(n_138), .Y(n_294) );
BUFx2_ASAP7_75t_L g321 ( .A(n_138), .Y(n_321) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_171), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_139), .B(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_139), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_139), .A2(n_241), .B(n_248), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_139), .B(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_139), .A2(n_502), .B(n_508), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_139), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_140), .A2(n_228), .B(n_229), .Y(n_227) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_140), .Y(n_268) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g250 ( .A(n_141), .Y(n_250) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_142), .B(n_143), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_167), .Y(n_146) );
INVx5_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx3_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx1_ASAP7_75t_L g236 ( .A(n_150), .Y(n_236) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_152), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
AND2x2_ASAP7_75t_L g169 ( .A(n_152), .B(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx1_ASAP7_75t_L g232 ( .A(n_152), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .C(n_161), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_156), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_156), .B(n_485), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_156), .A2(n_159), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
INVx2_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_159), .B(n_274), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_159), .A2(n_214), .B(n_515), .C(n_516), .Y(n_514) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_160), .B(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g499 ( .A(n_162), .Y(n_499) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_164), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_164), .A2(n_178), .B(n_271), .C(n_272), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_164), .A2(n_178), .B(n_453), .C(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_164), .A2(n_178), .B(n_461), .C(n_462), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_164), .A2(n_178), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_164), .A2(n_178), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_164), .A2(n_178), .B(n_529), .C(n_530), .Y(n_528) );
INVx4_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g168 ( .A(n_165), .B(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_165), .B(n_169), .Y(n_243) );
BUFx2_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
INVx1_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
AND2x2_ASAP7_75t_L g261 ( .A(n_173), .B(n_206), .Y(n_261) );
INVx2_ASAP7_75t_L g277 ( .A(n_173), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_173), .B(n_205), .Y(n_286) );
AND2x2_ASAP7_75t_L g365 ( .A(n_173), .B(n_294), .Y(n_365) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_187), .Y(n_173) );
INVx2_ASAP7_75t_L g195 ( .A(n_178), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_183), .B(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g463 ( .A(n_184), .Y(n_463) );
INVx2_ASAP7_75t_L g476 ( .A(n_185), .Y(n_476) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx1_ASAP7_75t_L g486 ( .A(n_186), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_222), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_189), .B(n_292), .Y(n_330) );
INVx1_ASAP7_75t_L g418 ( .A(n_189), .Y(n_418) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_205), .Y(n_189) );
AND2x2_ASAP7_75t_L g276 ( .A(n_190), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g290 ( .A(n_190), .B(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_190), .Y(n_319) );
OR2x2_ASAP7_75t_L g351 ( .A(n_190), .B(n_293), .Y(n_351) );
AND2x2_ASAP7_75t_L g359 ( .A(n_190), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g392 ( .A(n_190), .B(n_361), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_190), .B(n_261), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_190), .B(n_321), .Y(n_417) );
AND2x2_ASAP7_75t_L g423 ( .A(n_190), .B(n_310), .Y(n_423) );
INVx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g283 ( .A(n_191), .Y(n_283) );
AND2x2_ASAP7_75t_L g313 ( .A(n_191), .B(n_293), .Y(n_313) );
AND2x2_ASAP7_75t_L g346 ( .A(n_191), .B(n_306), .Y(n_346) );
AND2x2_ASAP7_75t_L g366 ( .A(n_191), .B(n_206), .Y(n_366) );
AND2x2_ASAP7_75t_L g400 ( .A(n_191), .B(n_266), .Y(n_400) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_203), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_202), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .C(n_201), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_201), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp5_ASAP7_75t_L g473 ( .A1(n_198), .A2(n_474), .B(n_475), .C(n_476), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_198), .A2(n_476), .B(n_506), .C(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g218 ( .A(n_202), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_202), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_202), .A2(n_254), .B(n_255), .Y(n_253) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_202), .A2(n_459), .B(n_466), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_202), .A2(n_243), .B(n_512), .C(n_513), .Y(n_511) );
AND2x4_ASAP7_75t_L g306 ( .A(n_205), .B(n_277), .Y(n_306) );
AND2x2_ASAP7_75t_L g317 ( .A(n_205), .B(n_313), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_205), .B(n_293), .Y(n_356) );
INVx2_ASAP7_75t_L g371 ( .A(n_205), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_205), .B(n_305), .Y(n_394) );
AND2x2_ASAP7_75t_L g413 ( .A(n_205), .B(n_365), .Y(n_413) );
INVx5_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_206), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_206), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g361 ( .A(n_206), .B(n_277), .Y(n_361) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_210), .B(n_217), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_215), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_218), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_221), .A2(n_470), .B(n_477), .Y(n_469) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
AND2x2_ASAP7_75t_L g284 ( .A(n_224), .B(n_267), .Y(n_284) );
INVx1_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_225), .B(n_240), .Y(n_264) );
OR2x2_ASAP7_75t_L g297 ( .A(n_225), .B(n_267), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_225), .B(n_267), .Y(n_302) );
AND2x2_ASAP7_75t_L g329 ( .A(n_225), .B(n_266), .Y(n_329) );
AND2x2_ASAP7_75t_L g381 ( .A(n_225), .B(n_239), .Y(n_381) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_226), .B(n_251), .Y(n_289) );
AND2x2_ASAP7_75t_L g325 ( .A(n_226), .B(n_240), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_233), .B(n_234), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_234), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_237), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g315 ( .A(n_238), .B(n_297), .Y(n_315) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_251), .Y(n_238) );
OAI322xp33_ASAP7_75t_L g280 ( .A1(n_239), .A2(n_281), .A3(n_285), .B1(n_287), .B2(n_290), .C1(n_295), .C2(n_303), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_239), .B(n_266), .Y(n_288) );
OR2x2_ASAP7_75t_L g298 ( .A(n_239), .B(n_252), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_239), .B(n_252), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_239), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_239), .B(n_267), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_239), .B(n_396), .Y(n_395) );
INVx5_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_240), .B(n_284), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_244), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_243), .A2(n_471), .B(n_472), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_243), .A2(n_503), .B(n_504), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g526 ( .A(n_250), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_251), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_251), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g340 ( .A(n_251), .B(n_267), .Y(n_340) );
AOI211xp5_ASAP7_75t_SL g368 ( .A1(n_251), .A2(n_369), .B(n_372), .C(n_384), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_251), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g406 ( .A(n_251), .B(n_381), .Y(n_406) );
INVx5_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g334 ( .A(n_252), .B(n_267), .Y(n_334) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
AND2x2_ASAP7_75t_L g383 ( .A(n_252), .B(n_381), .Y(n_383) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_252), .B(n_284), .Y(n_414) );
AND2x2_ASAP7_75t_L g421 ( .A(n_252), .B(n_380), .Y(n_421) );
OR2x6_ASAP7_75t_L g252 ( .A(n_253), .B(n_259), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B1(n_276), .B2(n_278), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_261), .B(n_283), .Y(n_331) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
OR2x2_ASAP7_75t_L g339 ( .A(n_264), .B(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_SL g387 ( .A1(n_264), .A2(n_388), .B1(n_390), .B2(n_391), .C(n_393), .Y(n_387) );
INVx2_ASAP7_75t_L g326 ( .A(n_265), .Y(n_326) );
AND2x2_ASAP7_75t_L g299 ( .A(n_266), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_266), .B(n_381), .Y(n_402) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g344 ( .A(n_267), .Y(n_344) );
AND2x2_ASAP7_75t_L g380 ( .A(n_267), .B(n_381), .Y(n_380) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_275), .Y(n_267) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_268), .A2(n_451), .B(n_457), .Y(n_450) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_268), .A2(n_480), .B(n_487), .Y(n_479) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_268), .A2(n_493), .B(n_500), .Y(n_492) );
AND2x2_ASAP7_75t_L g382 ( .A(n_276), .B(n_321), .Y(n_382) );
AND2x2_ASAP7_75t_L g292 ( .A(n_277), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_277), .B(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_279), .B(n_326), .Y(n_363) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g369 ( .A(n_282), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OR2x2_ASAP7_75t_L g355 ( .A(n_283), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g420 ( .A(n_283), .B(n_365), .Y(n_420) );
INVx2_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
NAND4xp25_ASAP7_75t_SL g416 ( .A(n_285), .B(n_417), .C(n_418), .D(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_286), .B(n_350), .Y(n_385) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_SL g422 ( .A(n_289), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_SL g384 ( .A1(n_290), .A2(n_353), .B(n_357), .C(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g379 ( .A(n_292), .B(n_371), .Y(n_379) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_293), .Y(n_305) );
INVx1_ASAP7_75t_L g360 ( .A(n_293), .Y(n_360) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B(n_299), .C(n_301), .Y(n_295) );
AND2x2_ASAP7_75t_L g316 ( .A(n_296), .B(n_300), .Y(n_316) );
OAI322xp33_ASAP7_75t_SL g354 ( .A1(n_296), .A2(n_355), .A3(n_357), .B1(n_358), .B2(n_362), .C1(n_363), .C2(n_364), .Y(n_354) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g376 ( .A(n_298), .B(n_302), .Y(n_376) );
INVx1_ASAP7_75t_L g357 ( .A(n_300), .Y(n_357) );
INVx1_ASAP7_75t_SL g375 ( .A(n_302), .Y(n_375) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_314), .B1(n_316), .B2(n_317), .C1(n_318), .C2(n_725), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_309), .B(n_311), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g397 ( .A1(n_309), .A2(n_371), .A3(n_376), .B1(n_398), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_324), .B1(n_348), .B2(n_352), .C(n_354), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
OAI222xp33_ASAP7_75t_L g327 ( .A1(n_315), .A2(n_328), .B1(n_330), .B2(n_331), .C1(n_332), .C2(n_335), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_317), .A2(n_324), .B1(n_394), .B2(n_395), .Y(n_393) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AOI211xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_327), .C(n_338), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g403 ( .A1(n_324), .A2(n_361), .B(n_404), .C(n_407), .Y(n_403) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_325), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g396 ( .A(n_329), .Y(n_396) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_336), .B(n_361), .Y(n_390) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_345), .Y(n_338) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_339), .A2(n_408), .B1(n_409), .B2(n_410), .C(n_411), .Y(n_407) );
INVxp33_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_343), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_350), .B(n_361), .Y(n_401) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_371), .Y(n_412) );
AND4x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_386), .C(n_403), .D(n_415), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B1(n_376), .B2(n_377), .C(n_378), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_382), .B2(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
INVx1_ASAP7_75t_SL g398 ( .A(n_383), .Y(n_398) );
NOR2xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_397), .Y(n_386) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_399), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_406), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g433 ( .A(n_428), .Y(n_433) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_429), .B(n_443), .Y(n_717) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g442 ( .A(n_430), .B(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_432), .A2(n_435), .B(n_722), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_441), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx6_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g720 ( .A(n_442), .Y(n_720) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g721 ( .A(n_445), .Y(n_721) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_631), .Y(n_445) );
NOR4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_573), .C(n_603), .D(n_613), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_488), .B(n_536), .C(n_563), .Y(n_447) );
OAI222xp33_ASAP7_75t_L g658 ( .A1(n_448), .A2(n_578), .B1(n_659), .B2(n_660), .C1(n_661), .C2(n_662), .Y(n_658) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_467), .Y(n_448) );
AOI33xp33_ASAP7_75t_L g584 ( .A1(n_449), .A2(n_571), .A3(n_572), .B1(n_585), .B2(n_590), .B3(n_592), .Y(n_584) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_449), .A2(n_642), .B(n_644), .C(n_646), .Y(n_641) );
OR2x2_ASAP7_75t_L g657 ( .A(n_449), .B(n_643), .Y(n_657) );
INVx1_ASAP7_75t_L g690 ( .A(n_449), .Y(n_690) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .Y(n_449) );
INVx2_ASAP7_75t_L g567 ( .A(n_450), .Y(n_567) );
AND2x2_ASAP7_75t_L g583 ( .A(n_450), .B(n_479), .Y(n_583) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_450), .Y(n_618) );
AND2x2_ASAP7_75t_L g647 ( .A(n_450), .B(n_458), .Y(n_647) );
INVx2_ASAP7_75t_L g547 ( .A(n_458), .Y(n_547) );
BUFx3_ASAP7_75t_L g555 ( .A(n_458), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_458), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g566 ( .A(n_458), .B(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_458), .B(n_468), .Y(n_595) );
AND2x2_ASAP7_75t_L g664 ( .A(n_458), .B(n_598), .Y(n_664) );
INVx2_ASAP7_75t_SL g558 ( .A(n_467), .Y(n_558) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_468), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g600 ( .A(n_468), .Y(n_600) );
AND2x2_ASAP7_75t_L g611 ( .A(n_468), .B(n_567), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_468), .B(n_596), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_468), .B(n_598), .Y(n_643) );
AND2x2_ASAP7_75t_L g702 ( .A(n_468), .B(n_647), .Y(n_702) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g572 ( .A(n_469), .B(n_479), .Y(n_572) );
AND2x2_ASAP7_75t_L g582 ( .A(n_469), .B(n_583), .Y(n_582) );
BUFx3_ASAP7_75t_L g604 ( .A(n_469), .Y(n_604) );
AND3x2_ASAP7_75t_L g663 ( .A(n_469), .B(n_664), .C(n_665), .Y(n_663) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_479), .Y(n_554) );
INVx1_ASAP7_75t_SL g598 ( .A(n_479), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_479), .B(n_547), .C(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_519), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_489), .A2(n_582), .B(n_634), .C(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_491), .B(n_510), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_491), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_SL g650 ( .A(n_491), .Y(n_650) );
AND2x2_ASAP7_75t_L g671 ( .A(n_491), .B(n_521), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_491), .B(n_580), .Y(n_699) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
AND2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_535), .Y(n_544) );
INVx2_ASAP7_75t_L g551 ( .A(n_492), .Y(n_551) );
AND2x2_ASAP7_75t_L g571 ( .A(n_492), .B(n_521), .Y(n_571) );
AND2x2_ASAP7_75t_L g621 ( .A(n_492), .B(n_510), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_492), .Y(n_625) );
INVx2_ASAP7_75t_SL g535 ( .A(n_501), .Y(n_535) );
BUFx2_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
AND2x2_ASAP7_75t_L g688 ( .A(n_501), .B(n_510), .Y(n_688) );
INVx3_ASAP7_75t_SL g521 ( .A(n_510), .Y(n_521) );
AND2x2_ASAP7_75t_L g543 ( .A(n_510), .B(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g550 ( .A(n_510), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g580 ( .A(n_510), .B(n_540), .Y(n_580) );
OR2x2_ASAP7_75t_L g589 ( .A(n_510), .B(n_535), .Y(n_589) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_510), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_510), .B(n_565), .Y(n_612) );
AND2x2_ASAP7_75t_L g640 ( .A(n_510), .B(n_523), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_510), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g678 ( .A(n_510), .B(n_522), .Y(n_678) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AND2x2_ASAP7_75t_L g602 ( .A(n_521), .B(n_551), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_521), .B(n_544), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_521), .B(n_565), .Y(n_648) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_535), .Y(n_522) );
AND2x2_ASAP7_75t_L g549 ( .A(n_523), .B(n_535), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_523), .B(n_578), .Y(n_577) );
BUFx3_ASAP7_75t_L g587 ( .A(n_523), .Y(n_587) );
OR2x2_ASAP7_75t_L g635 ( .A(n_523), .B(n_555), .Y(n_635) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_527), .B(n_534), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_525), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g541 ( .A(n_527), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_534), .Y(n_542) );
AND2x2_ASAP7_75t_L g570 ( .A(n_535), .B(n_540), .Y(n_570) );
INVx1_ASAP7_75t_L g578 ( .A(n_535), .Y(n_578) );
AND2x2_ASAP7_75t_L g673 ( .A(n_535), .B(n_551), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_545), .B1(n_548), .B2(n_552), .C1(n_556), .C2(n_559), .Y(n_536) );
INVx1_ASAP7_75t_L g668 ( .A(n_537), .Y(n_668) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
AND2x2_ASAP7_75t_L g564 ( .A(n_538), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g575 ( .A(n_538), .B(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_538), .B(n_566), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g613 ( .A1(n_538), .A2(n_614), .B1(n_619), .B2(n_620), .C1(n_628), .C2(n_630), .Y(n_613) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_540), .B(n_621), .Y(n_661) );
AND2x2_ASAP7_75t_L g672 ( .A(n_540), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g680 ( .A(n_543), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_545), .B(n_596), .Y(n_659) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_547), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_547), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx3_ASAP7_75t_L g562 ( .A(n_550), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_550), .A2(n_653), .B(n_656), .C(n_658), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_550), .B(n_587), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_550), .B(n_570), .Y(n_692) );
AND2x2_ASAP7_75t_L g565 ( .A(n_551), .B(n_561), .Y(n_565) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g592 ( .A(n_554), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_555), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g644 ( .A(n_555), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_583), .Y(n_683) );
INVx1_ASAP7_75t_L g695 ( .A(n_555), .Y(n_695) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_558), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g676 ( .A(n_561), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_566), .B(n_568), .C(n_572), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_564), .A2(n_594), .B1(n_609), .B2(n_612), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_565), .B(n_579), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_565), .B(n_587), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_566), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g629 ( .A(n_566), .Y(n_629) );
AND2x2_ASAP7_75t_L g636 ( .A(n_566), .B(n_616), .Y(n_636) );
INVx2_ASAP7_75t_L g597 ( .A(n_567), .Y(n_597) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NOR4xp25_ASAP7_75t_L g574 ( .A(n_571), .B(n_575), .C(n_576), .D(n_579), .Y(n_574) );
INVx1_ASAP7_75t_SL g645 ( .A(n_572), .Y(n_645) );
AND2x2_ASAP7_75t_L g689 ( .A(n_572), .B(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_581), .B(n_584), .C(n_593), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_580), .B(n_650), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_582), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
INVx1_ASAP7_75t_SL g655 ( .A(n_583), .Y(n_655) );
AND2x2_ASAP7_75t_L g694 ( .A(n_583), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_587), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_591), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_592), .B(n_617), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_599), .B(n_601), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g669 ( .A(n_596), .Y(n_669) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_L g697 ( .A(n_597), .Y(n_697) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_608), .Y(n_603) );
CKINVDCx16_ASAP7_75t_R g616 ( .A(n_604), .Y(n_616) );
OR2x2_ASAP7_75t_L g654 ( .A(n_604), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI21xp33_ASAP7_75t_SL g649 ( .A1(n_607), .A2(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_638), .B1(n_641), .B2(n_648), .C(n_649), .Y(n_637) );
INVx1_ASAP7_75t_SL g681 ( .A(n_612), .Y(n_681) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
OR2x2_ASAP7_75t_L g628 ( .A(n_616), .B(n_629), .Y(n_628) );
INVxp67_ASAP7_75t_L g665 ( .A(n_618), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_625), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g660 ( .A(n_621), .Y(n_660) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_624), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_666), .C(n_679), .D(n_691), .Y(n_631) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_633), .B(n_637), .C(n_652), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_635), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_642), .B(n_647), .Y(n_651) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_654), .A2(n_680), .B1(n_681), .B2(n_682), .C(n_684), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_656), .A2(n_671), .B(n_672), .C(n_674), .Y(n_670) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_657), .A2(n_675), .B1(n_677), .B2(n_678), .Y(n_674) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B(n_669), .C(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g685 ( .A(n_678), .Y(n_685) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_686), .B(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_693), .B1(n_696), .B2(n_698), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx3_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
endmodule