module fake_jpeg_29468_n_375 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_47),
.Y(n_135)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_68),
.Y(n_95)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_6),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_69),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_6),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_41),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_44),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_90),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_22),
.B(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_22),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_30),
.B(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_10),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_99),
.B(n_105),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_25),
.B1(n_17),
.B2(n_30),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_107),
.B1(n_84),
.B2(n_83),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_28),
.B1(n_37),
.B2(n_19),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_32),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_119),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_37),
.B1(n_11),
.B2(n_13),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_76),
.B1(n_74),
.B2(n_72),
.Y(n_156)
);

AND2x4_ASAP7_75t_SL g127 ( 
.A(n_54),
.B(n_25),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_52),
.B(n_25),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_137),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_55),
.B(n_5),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_1),
.Y(n_164)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_62),
.B1(n_84),
.B2(n_79),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_150),
.A2(n_179),
.B(n_157),
.C(n_172),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_95),
.B(n_58),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_154),
.A2(n_156),
.B1(n_160),
.B2(n_172),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_17),
.B(n_66),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_161),
.B(n_186),
.Y(n_212)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_169),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_168),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_187),
.Y(n_194)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_103),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_100),
.A2(n_107),
.B1(n_114),
.B2(n_113),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_143),
.B1(n_111),
.B2(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_177),
.B1(n_104),
.B2(n_115),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_142),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_111),
.A2(n_121),
.B1(n_109),
.B2(n_143),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_146),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_127),
.A2(n_145),
.B(n_92),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_93),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_136),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_129),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_130),
.B1(n_138),
.B2(n_97),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_170),
.B1(n_182),
.B2(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_104),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_220),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_104),
.A3(n_132),
.B1(n_97),
.B2(n_115),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_174),
.B1(n_184),
.B2(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_149),
.Y(n_208)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_150),
.B(n_186),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_178),
.B(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_159),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_152),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_153),
.B(n_151),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_226),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_197),
.B(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_231),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_230),
.B(n_253),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_161),
.B1(n_156),
.B2(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_161),
.B1(n_191),
.B2(n_162),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_222),
.A2(n_147),
.B1(n_158),
.B2(n_148),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_180),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_246),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_219),
.B(n_203),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_243),
.C(n_209),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_191),
.B1(n_170),
.B2(n_177),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_206),
.B1(n_205),
.B2(n_218),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_165),
.B(n_189),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_216),
.B(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_163),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_247),
.A2(n_193),
.B1(n_195),
.B2(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_202),
.A2(n_223),
.B1(n_199),
.B2(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_213),
.B(n_198),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_204),
.C(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_199),
.B(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_199),
.B(n_192),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_192),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_215),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_217),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_265),
.Y(n_283)
);

CKINVDCx10_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

NAND4xp25_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_271),
.C(n_244),
.D(n_240),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_254),
.B1(n_246),
.B2(n_247),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_204),
.C(n_211),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_224),
.C(n_221),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_216),
.B1(n_201),
.B2(n_195),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_277),
.B1(n_241),
.B2(n_236),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_229),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_280),
.A2(n_282),
.B1(n_296),
.B2(n_256),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_249),
.B1(n_234),
.B2(n_237),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_292),
.B1(n_294),
.B2(n_260),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_262),
.C(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_297),
.C(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_235),
.B1(n_233),
.B2(n_228),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_259),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_235),
.B1(n_233),
.B2(n_239),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_267),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_238),
.B1(n_252),
.B2(n_242),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_229),
.C(n_245),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_201),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_248),
.C(n_251),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_302),
.A2(n_282),
.B1(n_296),
.B2(n_280),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_274),
.B(n_267),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_304),
.A2(n_277),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_259),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_270),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_256),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_270),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_316),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_274),
.C(n_264),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_312),
.C(n_317),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_288),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_193),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_201),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_331),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_298),
.B(n_284),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_321),
.A2(n_304),
.B(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_295),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_325),
.C(n_333),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_302),
.A2(n_299),
.B1(n_291),
.B2(n_286),
.Y(n_327)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_315),
.B1(n_301),
.B2(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_336),
.B(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_322),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_343),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_305),
.C(n_308),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_333),
.C(n_328),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_332),
.B(n_310),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_346),
.B(n_349),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_337),
.A2(n_339),
.B(n_321),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_335),
.B(n_326),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_334),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_325),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_353),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_329),
.B(n_310),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_347),
.B(n_340),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_341),
.Y(n_358)
);

AO21x1_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_360),
.B(n_345),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_327),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_356),
.C(n_360),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_351),
.A2(n_334),
.B1(n_319),
.B2(n_338),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_361),
.B(n_348),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_357),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_365),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_364),
.B(n_366),
.Y(n_369)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_362),
.A2(n_358),
.B(n_348),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_368),
.B(n_367),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_369),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_371),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_342),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_343),
.B(n_345),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_331),
.Y(n_375)
);


endmodule