module fake_netlist_5_793_n_1775 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1775);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1775;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_24),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx11_ASAP7_75t_R g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_43),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_40),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_9),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_30),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_52),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_74),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_77),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_12),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_51),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_5),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_120),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_69),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_14),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_81),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_22),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_12),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_96),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_68),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_57),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_83),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_70),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_36),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_67),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_23),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_19),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_44),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_60),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_41),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_14),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_28),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_84),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_30),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_55),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_45),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_92),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_75),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_31),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_132),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_47),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_0),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_47),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_121),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_95),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_140),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_20),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_21),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_146),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_41),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_101),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_105),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_115),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_56),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_125),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_82),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_109),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_93),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_46),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_128),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_72),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_80),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_116),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_34),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_62),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_98),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_88),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_39),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_119),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_1),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_38),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_145),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_49),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_138),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_197),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_166),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_174),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_199),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_174),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_174),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_156),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_157),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_174),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_263),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_210),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_174),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_293),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_216),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_199),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_158),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_216),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_159),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_216),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_216),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_180),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_216),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_169),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_171),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_220),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_246),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_179),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_220),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_181),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_187),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_187),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_184),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_211),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_211),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_219),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_219),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_222),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_186),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_160),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_189),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_222),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_223),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_223),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_198),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_234),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_240),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_240),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_245),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_249),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_249),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_254),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_254),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_291),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_192),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_195),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_262),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_209),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_314),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_317),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_320),
.B(n_209),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_322),
.B(n_243),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_327),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_333),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_335),
.B(n_336),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_331),
.A2(n_161),
.B(n_155),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_349),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_309),
.B(n_198),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_355),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_309),
.B(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

NOR2x1_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_243),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_358),
.B(n_306),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_307),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_313),
.B(n_306),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_313),
.B(n_201),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_326),
.B(n_155),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_359),
.B(n_161),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_325),
.A2(n_246),
.B1(n_170),
.B2(n_206),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_326),
.B(n_204),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_360),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_323),
.A2(n_214),
.B1(n_256),
.B2(n_227),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_326),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_376),
.B(n_162),
.Y(n_444)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_321),
.B(n_162),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_371),
.B(n_208),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_341),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_341),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_320),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_339),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_376),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_411),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_212),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_407),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_434),
.A2(n_284),
.B1(n_267),
.B2(n_242),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_215),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_433),
.B(n_332),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

INVx8_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_442),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_345),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_377),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_418),
.B(n_217),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_445),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_445),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_413),
.B(n_316),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_418),
.B(n_308),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g481 ( 
.A1(n_404),
.A2(n_165),
.B(n_164),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_378),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_420),
.B(n_164),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_403),
.B(n_312),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_418),
.B(n_210),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_445),
.A2(n_200),
.B1(n_247),
.B2(n_255),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_406),
.B(n_316),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_407),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_434),
.A2(n_253),
.B1(n_173),
.B2(n_172),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_396),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_398),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_386),
.B(n_210),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_429),
.B(n_218),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_407),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_416),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_429),
.B(n_221),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_413),
.B(n_329),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

NOR2x1p5_ASAP7_75t_L g520 ( 
.A(n_402),
.B(n_232),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_390),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_440),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_426),
.B(n_346),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

AO22x1_ASAP7_75t_L g529 ( 
.A1(n_431),
.A2(n_351),
.B1(n_329),
.B2(n_372),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_438),
.B(n_210),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_420),
.B(n_226),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_449),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_393),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_409),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_436),
.B(n_228),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_407),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_390),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_390),
.Y(n_543)
);

INVxp33_ASAP7_75t_L g544 ( 
.A(n_441),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_387),
.B(n_229),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_441),
.A2(n_251),
.B1(n_175),
.B2(n_176),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_442),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_410),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_415),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_383),
.A2(n_370),
.B1(n_352),
.B2(n_351),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

AO22x2_ASAP7_75t_L g555 ( 
.A1(n_383),
.A2(n_296),
.B1(n_272),
.B2(n_273),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_431),
.B(n_348),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_383),
.B(n_238),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_383),
.B(n_244),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_419),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_431),
.A2(n_167),
.B(n_165),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_449),
.B(n_248),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_392),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_431),
.B(n_348),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_445),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_408),
.B(n_252),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_423),
.B(n_352),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_450),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_423),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_423),
.B(n_167),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_422),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_423),
.B(n_346),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_427),
.B(n_370),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_408),
.B(n_257),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_408),
.B(n_259),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_404),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_427),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_390),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_430),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_430),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_408),
.B(n_264),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_444),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_432),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_437),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_444),
.B(n_269),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_428),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_437),
.B(n_270),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_439),
.B(n_271),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_439),
.A2(n_247),
.B1(n_182),
.B2(n_177),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_390),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_443),
.B(n_274),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_499),
.B(n_485),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_574),
.B(n_444),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_468),
.B(n_310),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_462),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_556),
.B(n_444),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_569),
.A2(n_235),
.B1(n_279),
.B2(n_282),
.Y(n_607)
);

A2O1A1Ixp33_ASAP7_75t_L g608 ( 
.A1(n_578),
.A2(n_372),
.B(n_273),
.C(n_276),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_590),
.B(n_599),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_556),
.B(n_444),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_444),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_568),
.B(n_435),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_482),
.B(n_443),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_522),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_462),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_526),
.B(n_362),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_571),
.B(n_435),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_464),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_523),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_469),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_466),
.B(n_250),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_569),
.A2(n_285),
.B1(n_300),
.B2(n_294),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_590),
.B(n_250),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_576),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_590),
.B(n_250),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_590),
.B(n_250),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_516),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_530),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_473),
.B(n_178),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_435),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_514),
.B(n_435),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_517),
.B(n_435),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_480),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_538),
.B(n_435),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_535),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_537),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_477),
.B(n_362),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_547),
.B(n_447),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_537),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_466),
.B(n_250),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_466),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_541),
.B(n_447),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_461),
.B(n_185),
.Y(n_650)
);

INVx4_ASAP7_75t_SL g651 ( 
.A(n_484),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_447),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_549),
.B(n_447),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_597),
.A2(n_373),
.B(n_286),
.C(n_296),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_563),
.A2(n_404),
.B1(n_168),
.B2(n_190),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_590),
.B(n_250),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_549),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_480),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_467),
.B(n_168),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_492),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_560),
.A2(n_193),
.B1(n_279),
.B2(n_190),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_550),
.B(n_447),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_557),
.B(n_404),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_457),
.A2(n_200),
.B1(n_193),
.B2(n_182),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_492),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_561),
.B(n_399),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_561),
.B(n_399),
.Y(n_667)
);

BUFx5_ASAP7_75t_L g668 ( 
.A(n_599),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_493),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_551),
.B(n_188),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_590),
.B(n_250),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_599),
.B(n_250),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_551),
.B(n_194),
.Y(n_673)
);

AND2x6_ASAP7_75t_SL g674 ( 
.A(n_575),
.B(n_276),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_466),
.B(n_177),
.Y(n_675)
);

AO221x1_ASAP7_75t_L g676 ( 
.A1(n_501),
.A2(n_555),
.B1(n_286),
.B2(n_305),
.C(n_235),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_399),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_564),
.B(n_399),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_493),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_563),
.A2(n_297),
.B1(n_255),
.B2(n_258),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_599),
.B(n_494),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_567),
.B(n_399),
.Y(n_682)
);

NOR2x1p5_ASAP7_75t_L g683 ( 
.A(n_527),
.B(n_232),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_498),
.Y(n_684)
);

BUFx6f_ASAP7_75t_SL g685 ( 
.A(n_573),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_567),
.B(n_584),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_527),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_584),
.B(n_401),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_586),
.B(n_401),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_477),
.Y(n_690)
);

INVxp33_ASAP7_75t_SL g691 ( 
.A(n_576),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_498),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_563),
.A2(n_301),
.B1(n_265),
.B2(n_282),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_196),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_534),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_518),
.B(n_373),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_586),
.B(n_401),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_587),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_587),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_494),
.B(n_392),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_545),
.B(n_202),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_588),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_503),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_588),
.B(n_401),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_583),
.B(n_392),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_591),
.B(n_592),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_583),
.B(n_392),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_401),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_203),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_592),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_577),
.B(n_513),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_503),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_534),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_507),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_532),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_507),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_508),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_508),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_512),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_529),
.B(n_258),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_529),
.B(n_265),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_512),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_521),
.B(n_295),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_521),
.B(n_295),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_577),
.B(n_205),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_552),
.B(n_392),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_452),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_466),
.B(n_392),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_544),
.B(n_207),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_471),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_470),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_455),
.B(n_297),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_565),
.B(n_213),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_460),
.B(n_301),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_484),
.A2(n_305),
.B1(n_425),
.B2(n_417),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_546),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_533),
.B(n_224),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_474),
.B(n_417),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_471),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_597),
.A2(n_366),
.B(n_365),
.C(n_367),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_452),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_595),
.B(n_225),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_596),
.B(n_230),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_457),
.B(n_303),
.C(n_233),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_SL g745 ( 
.A1(n_475),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_554),
.B(n_277),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_456),
.B(n_417),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_554),
.B(n_287),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_456),
.B(n_425),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_500),
.B(n_425),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_573),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_453),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_453),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_500),
.B(n_448),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_458),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_454),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_600),
.B(n_239),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_515),
.B(n_448),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_472),
.Y(n_759)
);

INVx8_ASAP7_75t_L g760 ( 
.A(n_484),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_458),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_515),
.B(n_448),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_573),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_546),
.A2(n_381),
.B1(n_380),
.B2(n_379),
.C(n_375),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_454),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_484),
.A2(n_241),
.B1(n_266),
.B2(n_275),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_559),
.B(n_289),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_540),
.B(n_290),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_472),
.Y(n_769)
);

NAND2x1_ASAP7_75t_L g770 ( 
.A(n_648),
.B(n_490),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_632),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_602),
.B(n_559),
.Y(n_772)
);

BUFx4f_ASAP7_75t_L g773 ( 
.A(n_617),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_755),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_690),
.B(n_555),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_690),
.B(n_555),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_676),
.A2(n_555),
.B1(n_484),
.B2(n_575),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_610),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_615),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_620),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_605),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_636),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_614),
.B(n_484),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_755),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_606),
.B(n_540),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_641),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_629),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_644),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_605),
.Y(n_791)
);

BUFx12f_ASAP7_75t_SL g792 ( 
.A(n_643),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_616),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_687),
.B(n_475),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_696),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_713),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_634),
.B(n_484),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_711),
.A2(n_476),
.B1(n_475),
.B2(n_491),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_683),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_668),
.B(n_562),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_695),
.B(n_575),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_619),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_520),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_736),
.A2(n_476),
.B1(n_520),
.B2(n_593),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_479),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_SL g808 ( 
.A1(n_604),
.A2(n_763),
.B1(n_629),
.B2(n_691),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_755),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_657),
.B(n_575),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_698),
.B(n_575),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_668),
.B(n_562),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_619),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_680),
.A2(n_476),
.B1(n_536),
.B2(n_531),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_699),
.B(n_459),
.Y(n_815)
);

INVx5_ASAP7_75t_L g816 ( 
.A(n_760),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_668),
.B(n_581),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_642),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_621),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_702),
.B(n_459),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_621),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_755),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_622),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_729),
.B(n_570),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_611),
.B(n_581),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_691),
.Y(n_826)
);

OR2x2_ASAP7_75t_SL g827 ( 
.A(n_744),
.B(n_579),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_710),
.B(n_463),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_R g829 ( 
.A(n_763),
.B(n_481),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_623),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_715),
.B(n_580),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_670),
.B(n_589),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_623),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_673),
.B(n_278),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_761),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_650),
.B(n_280),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_764),
.B(n_283),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_714),
.B(n_463),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_668),
.B(n_648),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_639),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_718),
.B(n_465),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_658),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_668),
.B(n_582),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_751),
.B(n_365),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_668),
.B(n_582),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_668),
.B(n_594),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_725),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_760),
.B(n_366),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_648),
.B(n_594),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_719),
.B(n_465),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_686),
.B(n_706),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_612),
.A2(n_481),
.B1(n_572),
.B2(n_598),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_659),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_660),
.B(n_490),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_660),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_665),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_601),
.B(n_367),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_669),
.B(n_490),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_669),
.B(n_502),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_761),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_709),
.B(n_288),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_679),
.B(n_368),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_679),
.Y(n_866)
);

AND2x6_ASAP7_75t_SL g867 ( 
.A(n_701),
.B(n_368),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_684),
.B(n_502),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_608),
.A2(n_369),
.B(n_374),
.C(n_375),
.Y(n_869)
);

AND3x2_ASAP7_75t_SL g870 ( 
.A(n_664),
.B(n_1),
.C(n_3),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_684),
.B(n_502),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_733),
.B(n_369),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_692),
.B(n_572),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_692),
.B(n_572),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_663),
.B(n_495),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_703),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_659),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_703),
.B(n_598),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_712),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_712),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_716),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_655),
.A2(n_598),
.B1(n_304),
.B2(n_496),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_737),
.A2(n_585),
.B1(n_495),
.B2(n_504),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_716),
.B(n_478),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_717),
.Y(n_885)
);

BUFx6f_ASAP7_75t_SL g886 ( 
.A(n_659),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_717),
.B(n_478),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_722),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_720),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_722),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_761),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_727),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_741),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_760),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_741),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_752),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_721),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_613),
.B(n_495),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_753),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_608),
.B(n_374),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_734),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_705),
.A2(n_497),
.B1(n_483),
.B2(n_553),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_746),
.A2(n_585),
.B1(n_495),
.B2(n_504),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_753),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_756),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_732),
.B(n_292),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_685),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_705),
.B(n_298),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_765),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_765),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_760),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_685),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_723),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_707),
.A2(n_635),
.B(n_618),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_731),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_742),
.B(n_379),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_738),
.B(n_483),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_739),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_724),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_685),
.B(n_299),
.Y(n_922)
);

OR2x6_ASAP7_75t_SL g923 ( 
.A(n_607),
.B(n_380),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_759),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_746),
.Y(n_925)
);

AND2x6_ASAP7_75t_L g926 ( 
.A(n_603),
.B(n_495),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_769),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_693),
.B(n_486),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_707),
.B(n_486),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_654),
.B(n_381),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_666),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_681),
.A2(n_496),
.B1(n_497),
.B2(n_553),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_651),
.B(n_342),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_667),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_677),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_678),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_748),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_768),
.B(n_504),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_748),
.A2(n_585),
.B1(n_504),
.B2(n_509),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_682),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_688),
.Y(n_941)
);

NOR2x1p5_ASAP7_75t_L g942 ( 
.A(n_745),
.B(n_342),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_689),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_743),
.B(n_487),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_757),
.B(n_487),
.Y(n_945)
);

AND2x4_ASAP7_75t_SL g946 ( 
.A(n_625),
.B(n_504),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_697),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_704),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_767),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_SL g950 ( 
.A(n_661),
.B(n_343),
.C(n_347),
.Y(n_950)
);

OAI22xp33_ASAP7_75t_L g951 ( 
.A1(n_726),
.A2(n_681),
.B1(n_649),
.B2(n_652),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_645),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_651),
.B(n_343),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_726),
.A2(n_519),
.B1(n_488),
.B2(n_548),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_792),
.B(n_653),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_798),
.B(n_767),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_893),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_786),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_854),
.B(n_637),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_836),
.A2(n_675),
.B(n_624),
.C(n_647),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_836),
.B(n_638),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_893),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_797),
.B(n_773),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_797),
.B(n_766),
.Y(n_964)
);

CKINVDCx8_ASAP7_75t_R g965 ( 
.A(n_789),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_821),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_771),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_918),
.B(n_640),
.Y(n_968)
);

INVx3_ASAP7_75t_SL g969 ( 
.A(n_826),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_821),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_886),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_869),
.A2(n_740),
.B(n_662),
.C(n_708),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_864),
.B(n_747),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_902),
.B(n_872),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_786),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_869),
.A2(n_675),
.B(n_700),
.C(n_754),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_786),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_818),
.B(n_921),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_864),
.A2(n_647),
.B(n_624),
.C(n_672),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_795),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_917),
.A2(n_609),
.B(n_731),
.Y(n_981)
);

INVx5_ASAP7_75t_L g982 ( 
.A(n_895),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_832),
.A2(n_609),
.B1(n_735),
.B2(n_728),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_832),
.A2(n_672),
.B(n_758),
.C(n_750),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_846),
.B(n_834),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_824),
.B(n_651),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_818),
.B(n_749),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_SL g988 ( 
.A1(n_772),
.A2(n_630),
.B(n_627),
.C(n_671),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_896),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_876),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_917),
.A2(n_839),
.B(n_938),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_834),
.A2(n_762),
.B(n_631),
.C(n_671),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_917),
.A2(n_731),
.B(n_728),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_898),
.A2(n_519),
.B(n_548),
.C(n_488),
.Y(n_994)
);

CKINVDCx6p67_ASAP7_75t_R g995 ( 
.A(n_886),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_917),
.A2(n_731),
.B(n_470),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_876),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_805),
.B(n_731),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_L g999 ( 
.A1(n_775),
.A2(n_350),
.B1(n_354),
.B2(n_489),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_850),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_SL g1001 ( 
.A(n_816),
.B(n_656),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_898),
.A2(n_528),
.B(n_505),
.C(n_539),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_921),
.B(n_528),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_831),
.B(n_525),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_795),
.B(n_656),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_786),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_801),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_SL g1008 ( 
.A1(n_907),
.A2(n_489),
.B(n_505),
.C(n_506),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_860),
.B(n_631),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_889),
.B(n_4),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_906),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_860),
.B(n_506),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_SL g1013 ( 
.A1(n_899),
.A2(n_8),
.B(n_10),
.C(n_13),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_822),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_951),
.A2(n_510),
.B(n_511),
.C(n_531),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_837),
.A2(n_510),
.B(n_511),
.C(n_536),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_837),
.A2(n_539),
.B(n_543),
.C(n_542),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_877),
.A2(n_585),
.B1(n_509),
.B2(n_543),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_791),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_951),
.A2(n_8),
.B(n_13),
.C(n_15),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_793),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_831),
.B(n_585),
.C(n_543),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_907),
.A2(n_15),
.B(n_16),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_794),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_856),
.B(n_543),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_776),
.A2(n_509),
.B1(n_524),
.B2(n_525),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_802),
.A2(n_509),
.B(n_543),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_915),
.B(n_16),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_813),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_800),
.A2(n_542),
.B1(n_525),
.B2(n_524),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_839),
.A2(n_566),
.B(n_470),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_807),
.B(n_542),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_901),
.A2(n_509),
.B1(n_524),
.B2(n_525),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_906),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_822),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_930),
.A2(n_919),
.B(n_778),
.C(n_779),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_916),
.A2(n_566),
.B(n_470),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_910),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_780),
.B(n_524),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_781),
.B(n_524),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_909),
.A2(n_525),
.B(n_542),
.C(n_19),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_908),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_944),
.A2(n_542),
.B1(n_566),
.B2(n_63),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_803),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_802),
.A2(n_566),
.B(n_151),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_913),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_942),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_822),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_807),
.B(n_17),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_930),
.A2(n_18),
.B(n_23),
.C(n_25),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_811),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_822),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_783),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_782),
.B(n_25),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_812),
.A2(n_78),
.B(n_143),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_930),
.A2(n_27),
.B(n_29),
.C(n_31),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_819),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_812),
.A2(n_64),
.B(n_133),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_804),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_840),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_811),
.B(n_147),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_909),
.A2(n_27),
.B(n_29),
.C(n_32),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_823),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_925),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_796),
.A2(n_35),
.B(n_36),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_817),
.A2(n_86),
.B(n_114),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_830),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_784),
.B(n_37),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_840),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_788),
.B(n_37),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_817),
.A2(n_85),
.B(n_113),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_790),
.B(n_923),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_806),
.B(n_42),
.C(n_48),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_937),
.A2(n_42),
.B(n_49),
.C(n_50),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_865),
.B(n_53),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_945),
.A2(n_56),
.B(n_79),
.C(n_89),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_833),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_949),
.B(n_117),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_840),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_840),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_814),
.A2(n_94),
.B1(n_100),
.B2(n_108),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_841),
.A2(n_110),
.B(n_880),
.C(n_890),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_829),
.B(n_913),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_845),
.A2(n_849),
.B(n_848),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_891),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_810),
.B(n_950),
.C(n_777),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_814),
.A2(n_799),
.B1(n_816),
.B2(n_924),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_845),
.A2(n_848),
.B(n_849),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_842),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_774),
.B(n_835),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_858),
.A2(n_866),
.B(n_859),
.C(n_885),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_844),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_803),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_774),
.B(n_835),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_808),
.B(n_847),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_803),
.B(n_901),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_SL g1098 ( 
.A1(n_899),
.A2(n_888),
.B(n_873),
.C(n_861),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_985),
.A2(n_829),
.B1(n_953),
.B2(n_933),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1027),
.A2(n_855),
.B(n_852),
.Y(n_1100)
);

AO21x2_ASAP7_75t_L g1101 ( 
.A1(n_1017),
.A2(n_785),
.B(n_883),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_966),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1085),
.A2(n_852),
.B(n_770),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1004),
.A2(n_873),
.B(n_861),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1033),
.A2(n_827),
.B1(n_777),
.B2(n_924),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_961),
.A2(n_946),
.B(n_950),
.C(n_934),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_960),
.A2(n_816),
.B(n_928),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1089),
.A2(n_903),
.B(n_878),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_974),
.B(n_922),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1023),
.B(n_940),
.C(n_943),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_970),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_959),
.B(n_936),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_990),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_967),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_979),
.A2(n_929),
.B(n_932),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_968),
.A2(n_816),
.B(n_931),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_991),
.A2(n_874),
.B(n_857),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_1020),
.A2(n_935),
.B(n_941),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_978),
.B(n_980),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1088),
.A2(n_887),
.B(n_884),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1074),
.B(n_914),
.C(n_867),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_997),
.B(n_927),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_982),
.B(n_809),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_973),
.A2(n_947),
.B(n_948),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_973),
.A2(n_871),
.B(n_868),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1019),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1021),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1024),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1015),
.A2(n_862),
.B(n_932),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1003),
.B(n_881),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_992),
.A2(n_843),
.B(n_853),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1008),
.A2(n_904),
.B(n_939),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1029),
.Y(n_1133)
);

NAND2x1_ASAP7_75t_L g1134 ( 
.A(n_975),
.B(n_809),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1073),
.A2(n_870),
.B1(n_933),
.B2(n_879),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1063),
.B(n_838),
.C(n_815),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_984),
.A2(n_820),
.B(n_828),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_987),
.B(n_952),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1058),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1050),
.B(n_920),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1068),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1090),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1005),
.B(n_952),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_965),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_982),
.Y(n_1145)
);

AO32x2_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_882),
.A3(n_870),
.B1(n_825),
.B2(n_875),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1037),
.A2(n_895),
.B(n_912),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_895),
.B(n_912),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1054),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1005),
.B(n_1060),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_998),
.A2(n_911),
.B(n_894),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_977),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1082),
.A2(n_825),
.A3(n_875),
.B1(n_787),
.B2(n_954),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1045),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1052),
.B(n_900),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1064),
.B(n_952),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1015),
.A2(n_954),
.B(n_905),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1020),
.A2(n_892),
.B(n_897),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_988),
.A2(n_863),
.B(n_825),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_1042),
.A2(n_825),
.A3(n_875),
.B(n_787),
.Y(n_1160)
);

OAI22x1_ASAP7_75t_L g1161 ( 
.A1(n_1073),
.A2(n_863),
.B1(n_851),
.B2(n_825),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1078),
.B(n_952),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1026),
.A2(n_851),
.B(n_895),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1098),
.A2(n_787),
.B(n_875),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1093),
.B(n_891),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1012),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_976),
.A2(n_912),
.B(n_851),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1066),
.A2(n_891),
.B1(n_912),
.B2(n_787),
.C(n_926),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1092),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_976),
.A2(n_891),
.B(n_926),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_964),
.B(n_926),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_957),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1038),
.A2(n_926),
.B(n_1092),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_962),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1079),
.A2(n_926),
.B(n_1087),
.C(n_1010),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_963),
.B(n_955),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_994),
.A2(n_1002),
.B(n_1031),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_955),
.A2(n_1097),
.B1(n_1062),
.B2(n_1079),
.Y(n_1178)
);

BUFx8_ASAP7_75t_L g1179 ( 
.A(n_1047),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1009),
.B(n_989),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1011),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_986),
.A2(n_1065),
.B(n_1075),
.C(n_1026),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1034),
.B(n_1035),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1039),
.B(n_1052),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_SL g1185 ( 
.A(n_982),
.B(n_1049),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1022),
.A2(n_1016),
.B(n_1083),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_956),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_969),
.B(n_1096),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1083),
.A2(n_1006),
.B(n_1044),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1010),
.B(n_1028),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_971),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_981),
.A2(n_993),
.B(n_1033),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_994),
.A2(n_1002),
.B(n_972),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_972),
.A2(n_1046),
.B(n_1018),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1051),
.A2(n_1057),
.B1(n_1048),
.B2(n_1028),
.C(n_1071),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1040),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1076),
.B(n_1094),
.Y(n_1197)
);

AO21x1_ASAP7_75t_L g1198 ( 
.A1(n_1077),
.A2(n_999),
.B(n_1056),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1055),
.B(n_1069),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1006),
.A2(n_996),
.B(n_982),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1084),
.A2(n_1025),
.B(n_999),
.C(n_1001),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1007),
.B(n_1043),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1032),
.A2(n_1041),
.B(n_1072),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1080),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1086),
.B(n_958),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1086),
.A2(n_1036),
.B1(n_1049),
.B2(n_977),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_995),
.B(n_958),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_975),
.B(n_1061),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1059),
.A2(n_1067),
.B(n_1053),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1061),
.A2(n_1013),
.A3(n_1095),
.B(n_1091),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1014),
.A2(n_1070),
.B(n_1081),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_SL g1212 ( 
.A1(n_977),
.A2(n_1036),
.B(n_1049),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_977),
.A2(n_1036),
.B(n_1049),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1036),
.A2(n_1014),
.B(n_1081),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_971),
.B(n_1000),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_960),
.A2(n_648),
.B(n_959),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_960),
.A2(n_648),
.B(n_959),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_985),
.A2(n_602),
.B(n_836),
.Y(n_1218)
);

NOR2x1_ASAP7_75t_SL g1219 ( 
.A(n_982),
.B(n_816),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_974),
.B(n_516),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1027),
.A2(n_1089),
.B(n_1085),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_979),
.A2(n_602),
.B(n_960),
.Y(n_1222)
);

AO21x1_ASAP7_75t_L g1223 ( 
.A1(n_961),
.A2(n_602),
.B(n_1020),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_966),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1017),
.A2(n_1042),
.A3(n_960),
.B(n_961),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1074),
.A2(n_602),
.B1(n_832),
.B2(n_1073),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_966),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_L g1228 ( 
.A1(n_961),
.A2(n_602),
.B(n_836),
.C(n_864),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1033),
.A2(n_602),
.B1(n_960),
.B2(n_974),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_974),
.A2(n_602),
.B1(n_773),
.B2(n_526),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_980),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1094),
.B(n_1052),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1027),
.A2(n_1089),
.B(n_1085),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_979),
.A2(n_602),
.B(n_960),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_980),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_961),
.B(n_854),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_985),
.B(n_773),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_961),
.B(n_854),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1017),
.A2(n_1042),
.A3(n_960),
.B(n_961),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1141),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1231),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1237),
.B(n_1190),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1142),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1218),
.A2(n_1109),
.B1(n_1199),
.B2(n_1226),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1222),
.A2(n_1234),
.B(n_1217),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1235),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1114),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1228),
.A2(n_1110),
.B(n_1236),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1140),
.B(n_1166),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_1191),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1187),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_L g1252 ( 
.A(n_1188),
.B(n_1230),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1155),
.B(n_1176),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1238),
.B(n_1220),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1144),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1179),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1223),
.A2(n_1198),
.A3(n_1158),
.B(n_1168),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1195),
.B(n_1121),
.C(n_1175),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1234),
.A2(n_1135),
.B1(n_1229),
.B2(n_1105),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1229),
.A2(n_1105),
.B1(n_1112),
.B2(n_1169),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1197),
.B(n_1232),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1167),
.A2(n_1192),
.B(n_1170),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1143),
.Y(n_1263)
);

INVx4_ASAP7_75t_SL g1264 ( 
.A(n_1210),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1179),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1112),
.A2(n_1178),
.B1(n_1138),
.B2(n_1150),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1099),
.A2(n_1106),
.B1(n_1143),
.B2(n_1119),
.Y(n_1267)
);

AOI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_1171),
.B(n_1150),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1107),
.A2(n_1164),
.B(n_1186),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1207),
.B(n_1232),
.Y(n_1270)
);

CKINVDCx6p67_ASAP7_75t_R g1271 ( 
.A(n_1215),
.Y(n_1271)
);

AO21x2_ASAP7_75t_L g1272 ( 
.A1(n_1186),
.A2(n_1120),
.B(n_1189),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1154),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1126),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1122),
.B(n_1111),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1216),
.A2(n_1131),
.B(n_1137),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1152),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1124),
.A2(n_1116),
.B(n_1203),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1209),
.A2(n_1148),
.B(n_1103),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1202),
.B(n_1102),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1177),
.A2(n_1194),
.B(n_1100),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1108),
.A2(n_1147),
.B(n_1159),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1203),
.A2(n_1157),
.B(n_1151),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_L g1284 ( 
.A1(n_1182),
.A2(n_1118),
.B1(n_1227),
.B2(n_1113),
.C(n_1224),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1118),
.C(n_1115),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1180),
.B(n_1184),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1161),
.A2(n_1125),
.A3(n_1213),
.B(n_1163),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1129),
.A2(n_1104),
.B(n_1125),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1115),
.A2(n_1201),
.B(n_1130),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_SL g1291 ( 
.A1(n_1212),
.A2(n_1185),
.B(n_1214),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1127),
.A2(n_1139),
.B1(n_1133),
.B2(n_1128),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1215),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1200),
.A2(n_1211),
.B(n_1214),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1206),
.A2(n_1196),
.A3(n_1130),
.B(n_1153),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1206),
.A2(n_1156),
.B(n_1162),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1204),
.B(n_1172),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1146),
.A2(n_1153),
.B1(n_1219),
.B2(n_1149),
.Y(n_1298)
);

AO21x2_ASAP7_75t_L g1299 ( 
.A1(n_1132),
.A2(n_1101),
.B(n_1165),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1152),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1152),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1156),
.A2(n_1162),
.B(n_1165),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1174),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1123),
.A2(n_1183),
.B(n_1205),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1205),
.B(n_1181),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1183),
.A2(n_1146),
.B1(n_1123),
.B2(n_1208),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1208),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1134),
.A2(n_1101),
.B(n_1160),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1210),
.Y(n_1309)
);

OAI221xp5_ASAP7_75t_L g1310 ( 
.A1(n_1225),
.A2(n_602),
.B1(n_604),
.B2(n_836),
.C(n_864),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1210),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1160),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1225),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1239),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1239),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1228),
.B(n_602),
.C(n_836),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1145),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1163),
.B(n_1167),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1190),
.B(n_602),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1228),
.A2(n_602),
.B(n_836),
.Y(n_1320)
);

AOI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1228),
.A2(n_602),
.B(n_836),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1141),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1141),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1222),
.A2(n_960),
.B(n_1234),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1141),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1152),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1141),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1141),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1190),
.B(n_602),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1141),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_604),
.B2(n_836),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1222),
.A2(n_960),
.B(n_1234),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1141),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1222),
.A2(n_960),
.B(n_1234),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_1218),
.B2(n_1023),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_1218),
.B2(n_1023),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1221),
.A2(n_1233),
.B(n_1117),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1141),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1152),
.B(n_982),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1141),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1141),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_1218),
.B2(n_1023),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_SL g1343 ( 
.A(n_1228),
.B(n_602),
.C(n_1218),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_1238),
.B2(n_1236),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1141),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1166),
.B(n_1187),
.Y(n_1346)
);

BUFx2_ASAP7_75t_R g1347 ( 
.A(n_1144),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1228),
.A2(n_602),
.B(n_836),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1141),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1191),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1193),
.A2(n_1173),
.B(n_1222),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1190),
.A2(n_602),
.B1(n_604),
.B2(n_836),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1193),
.A2(n_1173),
.B(n_1222),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1114),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1222),
.A2(n_960),
.B(n_1234),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1191),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1114),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1141),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1175),
.A2(n_960),
.B(n_1063),
.C(n_979),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1143),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1222),
.A2(n_960),
.B(n_1234),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1152),
.B(n_982),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1228),
.B(n_602),
.C(n_836),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1255),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1247),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1331),
.A2(n_1352),
.B1(n_1319),
.B2(n_1329),
.Y(n_1366)
);

OA22x2_ASAP7_75t_L g1367 ( 
.A1(n_1244),
.A2(n_1348),
.B1(n_1320),
.B2(n_1251),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1276),
.A2(n_1310),
.B(n_1321),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1319),
.A2(n_1329),
.B1(n_1342),
.B2(n_1335),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1316),
.A2(n_1363),
.B(n_1362),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1346),
.B(n_1263),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1278),
.A2(n_1282),
.B(n_1289),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1274),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1339),
.A2(n_1362),
.B(n_1343),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1283),
.A2(n_1245),
.B(n_1248),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1301),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1247),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1263),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1360),
.B(n_1275),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1324),
.A2(n_1361),
.B(n_1334),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1261),
.B(n_1249),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1360),
.B(n_1286),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1255),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1332),
.A2(n_1355),
.B(n_1258),
.C(n_1342),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1280),
.B(n_1254),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1280),
.B(n_1270),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1359),
.A2(n_1318),
.B(n_1272),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1335),
.A2(n_1336),
.B1(n_1259),
.B2(n_1344),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1301),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_1250),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1359),
.A2(n_1318),
.B(n_1272),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1277),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1336),
.A2(n_1259),
.B1(n_1344),
.B2(n_1252),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1292),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_1241),
.B1(n_1246),
.B2(n_1318),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1356),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1270),
.B(n_1297),
.Y(n_1398)
);

INVxp33_ASAP7_75t_L g1399 ( 
.A(n_1273),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1339),
.A2(n_1343),
.B(n_1277),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1315),
.A2(n_1267),
.B1(n_1357),
.B2(n_1354),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1266),
.B(n_1323),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1266),
.A2(n_1285),
.B(n_1268),
.C(n_1305),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1337),
.A2(n_1311),
.B(n_1279),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1297),
.B(n_1325),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1284),
.A2(n_1298),
.B(n_1313),
.C(n_1358),
.Y(n_1406)
);

INVx3_ASAP7_75t_SL g1407 ( 
.A(n_1256),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1354),
.A2(n_1357),
.B1(n_1271),
.B2(n_1293),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1240),
.A2(n_1243),
.B1(n_1349),
.B2(n_1345),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1305),
.B(n_1330),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1262),
.A2(n_1285),
.B(n_1290),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1347),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1322),
.A2(n_1327),
.B(n_1340),
.C(n_1333),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1303),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1300),
.B(n_1296),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1277),
.B(n_1326),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1277),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1330),
.B(n_1341),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1328),
.A2(n_1338),
.B(n_1262),
.C(n_1291),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1295),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1295),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1308),
.A2(n_1294),
.B(n_1304),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1303),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1326),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1302),
.A2(n_1264),
.B(n_1257),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1295),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1326),
.A2(n_1307),
.B(n_1300),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1264),
.A2(n_1257),
.B(n_1269),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1356),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1306),
.A2(n_1290),
.B(n_1317),
.C(n_1288),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_R g1431 ( 
.A(n_1265),
.B(n_1307),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1265),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1287),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1290),
.B(n_1298),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1350),
.A2(n_1256),
.B1(n_1312),
.B2(n_1353),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1313),
.B(n_1257),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1257),
.B(n_1287),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1299),
.B(n_1309),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1312),
.B(n_1299),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1281),
.Y(n_1440)
);

BUFx8_ASAP7_75t_L g1441 ( 
.A(n_1351),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1281),
.B(n_1319),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1253),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1255),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1331),
.B(n_1352),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1331),
.A2(n_1352),
.B1(n_1319),
.B2(n_1329),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1331),
.A2(n_1352),
.B1(n_1319),
.B2(n_1329),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1331),
.A2(n_602),
.B(n_1228),
.C(n_1352),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1319),
.B(n_1329),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1314),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1319),
.B(n_1329),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1310),
.A2(n_602),
.B(n_1228),
.C(n_1319),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1441),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1368),
.A2(n_1411),
.B(n_1388),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1392),
.B(n_1381),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1421),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1450),
.A2(n_1454),
.B(n_1385),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1446),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1442),
.B(n_1426),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_1373),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1441),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1404),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1385),
.A2(n_1450),
.B(n_1430),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1452),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1415),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1415),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1425),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1375),
.B(n_1437),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1446),
.B(n_1366),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1375),
.B(n_1428),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1378),
.B(n_1395),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1438),
.A2(n_1436),
.B(n_1406),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1410),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1425),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1375),
.B(n_1428),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1428),
.B(n_1425),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1447),
.A2(n_1448),
.B1(n_1369),
.B2(n_1389),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1402),
.B(n_1380),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1419),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1418),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1371),
.B(n_1403),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1406),
.A2(n_1394),
.B(n_1370),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1372),
.A2(n_1422),
.B(n_1427),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1439),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1372),
.B(n_1405),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1435),
.B(n_1396),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1401),
.A2(n_1374),
.B(n_1409),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1397),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1413),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1367),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1367),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1386),
.B(n_1449),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1443),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1491),
.B(n_1445),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1491),
.B(n_1379),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1479),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1490),
.B(n_1399),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1482),
.A2(n_1391),
.B1(n_1397),
.B2(n_1408),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1491),
.B(n_1473),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1382),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1458),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1488),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1473),
.B(n_1398),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1462),
.B(n_1399),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1482),
.A2(n_1400),
.B1(n_1423),
.B2(n_1429),
.C(n_1414),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1387),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1459),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1469),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1463),
.B(n_1390),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1478),
.B(n_1417),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1460),
.A2(n_1429),
.B1(n_1432),
.B2(n_1414),
.C(n_1416),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1478),
.B(n_1393),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1475),
.B(n_1480),
.Y(n_1520)
);

OR2x2_ASAP7_75t_SL g1521 ( 
.A(n_1492),
.B(n_1496),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1465),
.B(n_1393),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1469),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1474),
.A2(n_1377),
.B1(n_1365),
.B2(n_1444),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1463),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1507),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1507),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1505),
.B(n_1465),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1504),
.A2(n_1460),
.B1(n_1497),
.B2(n_1486),
.C(n_1496),
.Y(n_1532)
);

NOR4xp25_ASAP7_75t_SL g1533 ( 
.A(n_1518),
.B(n_1416),
.C(n_1472),
.D(n_1495),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1507),
.Y(n_1534)
);

OAI33xp33_ASAP7_75t_L g1535 ( 
.A1(n_1525),
.A2(n_1486),
.A3(n_1497),
.B1(n_1483),
.B2(n_1495),
.B3(n_1489),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1526),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1504),
.A2(n_1497),
.B1(n_1496),
.B2(n_1468),
.C(n_1484),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1512),
.A2(n_1487),
.B1(n_1468),
.B2(n_1461),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1505),
.B(n_1466),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1518),
.A2(n_1487),
.B1(n_1461),
.B2(n_1468),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1512),
.B(n_1496),
.C(n_1495),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1509),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1502),
.B(n_1471),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1514),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1525),
.A2(n_1487),
.B1(n_1468),
.B2(n_1461),
.Y(n_1546)
);

OA222x2_ASAP7_75t_L g1547 ( 
.A1(n_1521),
.A2(n_1492),
.B1(n_1479),
.B2(n_1484),
.C1(n_1471),
.C2(n_1487),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1523),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1513),
.B(n_1489),
.C(n_1492),
.Y(n_1549)
);

OAI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1513),
.A2(n_1483),
.B(n_1456),
.C(n_1499),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1511),
.B(n_1499),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1502),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1516),
.A2(n_1487),
.B1(n_1468),
.B2(n_1461),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1502),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1432),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1516),
.A2(n_1461),
.B1(n_1477),
.B2(n_1493),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1466),
.Y(n_1558)
);

AOI211xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1508),
.A2(n_1457),
.B(n_1517),
.C(n_1519),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1516),
.A2(n_1461),
.B1(n_1477),
.B2(n_1493),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1500),
.A2(n_1457),
.B1(n_1498),
.B2(n_1476),
.C(n_1485),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1500),
.A2(n_1457),
.B1(n_1498),
.B2(n_1476),
.C(n_1485),
.Y(n_1562)
);

OAI31xp33_ASAP7_75t_L g1563 ( 
.A1(n_1503),
.A2(n_1457),
.A3(n_1455),
.B(n_1464),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1516),
.A2(n_1477),
.B1(n_1493),
.B2(n_1455),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1555),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1555),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1555),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1549),
.B(n_1455),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1527),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_SL g1571 ( 
.A(n_1533),
.B(n_1494),
.C(n_1503),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1531),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1528),
.Y(n_1575)
);

INVx4_ASAP7_75t_SL g1576 ( 
.A(n_1555),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1534),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1555),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1542),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1544),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1529),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1530),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1501),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1542),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1552),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1552),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1591)
);

INVx6_ASAP7_75t_L g1592 ( 
.A(n_1544),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1540),
.A2(n_1546),
.B(n_1538),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1545),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1529),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1532),
.B(n_1456),
.C(n_1376),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1529),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1543),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1535),
.A2(n_1493),
.B(n_1431),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1585),
.B(n_1584),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1570),
.Y(n_1603)
);

O2A1O1Ixp5_ASAP7_75t_SL g1604 ( 
.A1(n_1593),
.A2(n_1550),
.B(n_1515),
.C(n_1524),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1570),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1568),
.B(n_1501),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1572),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1544),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1494),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1522),
.Y(n_1612)
);

AOI33xp33_ASAP7_75t_L g1613 ( 
.A1(n_1586),
.A2(n_1564),
.A3(n_1560),
.B1(n_1557),
.B2(n_1537),
.B3(n_1533),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1521),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1596),
.B(n_1563),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1617)
);

AOI221x1_ASAP7_75t_L g1618 ( 
.A1(n_1571),
.A2(n_1541),
.B1(n_1515),
.B2(n_1524),
.C(n_1519),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1599),
.A2(n_1541),
.B(n_1553),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1536),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1575),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1520),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1576),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1589),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1575),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1592),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1592),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1565),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1586),
.B(n_1562),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1581),
.B(n_1521),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1574),
.B(n_1581),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_SL g1633 ( 
.A(n_1588),
.B(n_1464),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1579),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1574),
.B(n_1520),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1591),
.B(n_1506),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1565),
.B(n_1530),
.Y(n_1638)
);

NAND4xp25_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1563),
.C(n_1559),
.D(n_1457),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1588),
.B(n_1554),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1574),
.B(n_1567),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1579),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1642),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1506),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1623),
.Y(n_1645)
);

AOI322xp5_ASAP7_75t_L g1646 ( 
.A1(n_1630),
.A2(n_1505),
.A3(n_1520),
.B1(n_1558),
.B2(n_1548),
.C1(n_1506),
.C2(n_1574),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1510),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1609),
.B(n_1567),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1600),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1623),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1510),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1566),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1623),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1606),
.B(n_1510),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1624),
.B(n_1588),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1609),
.B(n_1588),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1641),
.B(n_1566),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1498),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1603),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1566),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1641),
.B(n_1578),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1601),
.B(n_1578),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1616),
.B(n_1578),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1578),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1605),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1608),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1610),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1616),
.B(n_1607),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1580),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1611),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1639),
.B(n_1407),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1615),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1621),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1618),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1645),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1657),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1670),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1650),
.B(n_1633),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1671),
.B(n_1629),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1648),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1648),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1672),
.B(n_1651),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1672),
.B(n_1628),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1658),
.Y(n_1691)
);

CKINVDCx16_ASAP7_75t_R g1692 ( 
.A(n_1674),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1650),
.B(n_1620),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1665),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1659),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1643),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1659),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1663),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1652),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1662),
.A2(n_1614),
.B1(n_1626),
.B2(n_1627),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1660),
.B(n_1407),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1652),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1645),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1682),
.A2(n_1700),
.B1(n_1701),
.B2(n_1686),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1691),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1707)
);

OAI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1679),
.A2(n_1644),
.B1(n_1657),
.B2(n_1656),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1692),
.A2(n_1658),
.B1(n_1676),
.B2(n_1663),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1695),
.B(n_1647),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1697),
.B(n_1666),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1694),
.B1(n_1684),
.B2(n_1653),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1685),
.A2(n_1664),
.B1(n_1667),
.B2(n_1653),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1681),
.A2(n_1655),
.B1(n_1645),
.B2(n_1640),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1693),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1718)
);

OAI322xp33_ASAP7_75t_L g1719 ( 
.A1(n_1690),
.A2(n_1677),
.A3(n_1668),
.B1(n_1661),
.B2(n_1678),
.C1(n_1669),
.C2(n_1649),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1681),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1693),
.A2(n_1604),
.B1(n_1667),
.B2(n_1464),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1717),
.Y(n_1723)
);

NOR2xp67_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1683),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1706),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1707),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1721),
.A2(n_1703),
.B1(n_1693),
.B2(n_1683),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1714),
.B(n_1703),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1705),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1722),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1711),
.B(n_1688),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1723),
.B(n_1718),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1729),
.A2(n_1721),
.B1(n_1708),
.B2(n_1719),
.C(n_1716),
.Y(n_1735)
);

AOI221x1_ASAP7_75t_L g1736 ( 
.A1(n_1725),
.A2(n_1720),
.B1(n_1712),
.B2(n_1699),
.C(n_1696),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1727),
.A2(n_1710),
.B1(n_1688),
.B2(n_1646),
.C(n_1689),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1726),
.B(n_1702),
.C(n_1678),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1733),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1728),
.A2(n_1731),
.B1(n_1730),
.B2(n_1732),
.C(n_1661),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1732),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1735),
.A2(n_1724),
.B1(n_1668),
.B2(n_1677),
.C(n_1689),
.Y(n_1743)
);

XNOR2xp5_ASAP7_75t_L g1744 ( 
.A(n_1742),
.B(n_1364),
.Y(n_1744)
);

OAI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1737),
.A2(n_1612),
.B(n_1622),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1738),
.A2(n_1364),
.B(n_1444),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1734),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1741),
.C(n_1744),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1740),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1747),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1746),
.Y(n_1751)
);

NAND2xp33_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1739),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1747),
.Y(n_1753)
);

OAI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1749),
.A2(n_1736),
.B(n_1612),
.Y(n_1754)
);

AOI21xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1748),
.A2(n_1384),
.B(n_1675),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1752),
.B(n_1384),
.C(n_1412),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1751),
.Y(n_1757)
);

NAND4xp75_ASAP7_75t_L g1758 ( 
.A(n_1750),
.B(n_1622),
.C(n_1625),
.D(n_1635),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1754),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1753),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1755),
.B(n_1675),
.C(n_1638),
.Y(n_1761)
);

AND3x1_ASAP7_75t_L g1762 ( 
.A(n_1759),
.B(n_1756),
.C(n_1758),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1762),
.B(n_1761),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1763),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1760),
.B1(n_1620),
.B2(n_1634),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1764),
.A2(n_1634),
.B1(n_1592),
.B2(n_1636),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1582),
.B(n_1376),
.Y(n_1768)
);

OAI22x1_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1582),
.B1(n_1587),
.B2(n_1594),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1769),
.B1(n_1582),
.B2(n_1598),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1771),
.B(n_1595),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1772),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1598),
.B1(n_1595),
.B2(n_1597),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1393),
.B(n_1424),
.C(n_1597),
.Y(n_1775)
);


endmodule