module fake_jpeg_5509_n_275 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_24),
.B1(n_21),
.B2(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_29),
.B1(n_28),
.B2(n_35),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_25),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g92 ( 
.A(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_49),
.C(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_52),
.B1(n_48),
.B2(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_51),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_52),
.B1(n_32),
.B2(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_81),
.B1(n_71),
.B2(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_35),
.A3(n_32),
.B1(n_42),
.B2(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_62),
.Y(n_112)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_101),
.B1(n_115),
.B2(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_99),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_93),
.Y(n_117)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_61),
.C(n_70),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_113),
.C(n_88),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_114),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_91),
.B1(n_81),
.B2(n_79),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_33),
.C(n_46),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_43),
.B1(n_72),
.B2(n_73),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_118),
.C(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_74),
.C(n_91),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_137),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_127),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_76),
.C(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_112),
.B1(n_105),
.B2(n_99),
.Y(n_141)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_135),
.B1(n_90),
.B2(n_31),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_33),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_136),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_114),
.Y(n_132)
);

NAND2xp67_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_51),
.B(n_33),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_33),
.C(n_31),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_27),
.B(n_23),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_109),
.B1(n_111),
.B2(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_141),
.B1(n_147),
.B2(n_150),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_127),
.B1(n_23),
.B2(n_30),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_112),
.B1(n_109),
.B2(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_117),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_90),
.B1(n_19),
.B2(n_25),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_31),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_30),
.C(n_23),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_120),
.B1(n_135),
.B2(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_159),
.B1(n_116),
.B2(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_122),
.B(n_31),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_164),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_160),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_174),
.C(n_176),
.Y(n_193)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_172),
.B1(n_157),
.B2(n_14),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_129),
.B1(n_132),
.B2(n_119),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_30),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_30),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_25),
.C(n_19),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_15),
.C(n_16),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_184),
.B(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_146),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_187),
.B(n_189),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_146),
.B1(n_158),
.B2(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_192),
.B1(n_195),
.B2(n_168),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_153),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_200),
.C(n_177),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_203),
.B(n_184),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_0),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_13),
.Y(n_202)
);

AOI31xp67_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_167),
.A3(n_166),
.B(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_206),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_209),
.B(n_6),
.Y(n_232)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_169),
.B(n_163),
.C(n_182),
.D(n_7),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_200),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_6),
.B1(n_10),
.B2(n_9),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_217),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_218),
.B(n_219),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_185),
.B1(n_193),
.B2(n_187),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_229),
.B1(n_0),
.B2(n_1),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_232),
.B(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_215),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_193),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_5),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_R g239 ( 
.A(n_233),
.B(n_215),
.C(n_7),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_208),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_238),
.C(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_214),
.B1(n_7),
.B2(n_8),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_225),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_245),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_221),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_255),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_254),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_9),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_8),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_1),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_260),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_9),
.B(n_10),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_12),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_12),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_270),
.B(n_264),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.B(n_4),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_267),
.B(n_3),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_3),
.Y(n_275)
);


endmodule