module fake_jpeg_23772_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx6_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_25),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_14),
.B1(n_29),
.B2(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_43),
.B1(n_14),
.B2(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_44),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_11),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_51),
.B1(n_42),
.B2(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_46),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_64),
.B1(n_56),
.B2(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AOI21x1_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_40),
.B(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.C(n_59),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_9),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_53),
.B1(n_49),
.B2(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_31),
.B1(n_1),
.B2(n_7),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_1),
.B(n_2),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_67),
.B1(n_8),
.B2(n_9),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_5),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_76),
.Y(n_78)
);


endmodule