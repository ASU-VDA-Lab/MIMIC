module fake_jpeg_214_n_684 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_684);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_684;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_61),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_11),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_85),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_80),
.Y(n_148)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_71),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_11),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_10),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_101),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

INVx11_ASAP7_75t_SL g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_42),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_43),
.B(n_10),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_103),
.B(n_104),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_119),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_12),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_18),
.Y(n_139)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_32),
.Y(n_123)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_21),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_50),
.Y(n_208)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_131),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_137),
.B(n_149),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_139),
.B(n_182),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_59),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_110),
.A2(n_27),
.B1(n_56),
.B2(n_54),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_158),
.A2(n_164),
.B1(n_176),
.B2(n_200),
.Y(n_244)
);

BUFx16f_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_63),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_163),
.B(n_168),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_84),
.A2(n_27),
.B1(n_56),
.B2(n_54),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_73),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_57),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_175),
.B(n_0),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_76),
.A2(n_33),
.B1(n_57),
.B2(n_48),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_76),
.B(n_23),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_75),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_81),
.B(n_23),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_194),
.B(n_208),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_87),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_111),
.A2(n_21),
.B1(n_50),
.B2(n_46),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_95),
.A2(n_57),
.B1(n_48),
.B2(n_58),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_203),
.A2(n_72),
.B1(n_116),
.B2(n_102),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_209),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_72),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_126),
.B(n_36),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_220),
.Y(n_280)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_88),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_94),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_98),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_34),
.Y(n_263)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_219),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_36),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_223),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_90),
.B(n_46),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_14),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_161),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_227),
.B(n_236),
.C(n_258),
.Y(n_348)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_230),
.Y(n_346)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_231),
.Y(n_360)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_232),
.Y(n_361)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_234),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_121),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_134),
.B(n_41),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_240),
.B(n_268),
.Y(n_311)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_157),
.A2(n_114),
.B1(n_41),
.B2(n_45),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_247),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_195),
.A2(n_187),
.B1(n_136),
.B2(n_132),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

CKINVDCx9p33_ASAP7_75t_R g249 ( 
.A(n_152),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_249),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_131),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_250),
.B(n_285),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_195),
.A2(n_57),
.B1(n_74),
.B2(n_112),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_136),
.A2(n_57),
.B1(n_119),
.B2(n_112),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_177),
.A2(n_118),
.B1(n_115),
.B2(n_125),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_152),
.Y(n_254)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_141),
.A2(n_119),
.B1(n_113),
.B2(n_108),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_262),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_179),
.B(n_102),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_176),
.A2(n_116),
.B1(n_45),
.B2(n_34),
.Y(n_262)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_264),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_290),
.Y(n_317)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_174),
.Y(n_266)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_266),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_28),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_145),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_284),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_157),
.B(n_28),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_273),
.B(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_169),
.Y(n_276)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_203),
.A2(n_24),
.B1(n_0),
.B2(n_2),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_181),
.B1(n_290),
.B2(n_289),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_24),
.Y(n_278)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_165),
.Y(n_281)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_144),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_282),
.A2(n_287),
.B1(n_221),
.B2(n_199),
.Y(n_358)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_159),
.B(n_13),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_207),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_295),
.Y(n_322)
);

OA22x2_ASAP7_75t_L g290 ( 
.A1(n_186),
.A2(n_14),
.B1(n_5),
.B2(n_9),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_148),
.B(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_291),
.B(n_292),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_148),
.B(n_5),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_156),
.Y(n_293)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_135),
.B(n_5),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_301),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_9),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_171),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_297),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_213),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_302),
.Y(n_329)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_220),
.B(n_13),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_167),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_178),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_307),
.Y(n_349)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_216),
.Y(n_369)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_236),
.B(n_142),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_308),
.B(n_358),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_153),
.C(n_162),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_314),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_150),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_310),
.B(n_328),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_SL g314 ( 
.A(n_265),
.B(n_138),
.C(n_198),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_235),
.B(n_143),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_316),
.B(n_332),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_248),
.B(n_140),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_320),
.B(n_216),
.CI(n_142),
.CON(n_416),
.SN(n_416)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_188),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_184),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_334),
.A2(n_337),
.B1(n_341),
.B2(n_289),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_277),
.A2(n_181),
.B1(n_218),
.B2(n_212),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_244),
.A2(n_237),
.B1(n_241),
.B2(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_246),
.B(n_199),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_365),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_251),
.A2(n_191),
.B(n_198),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_353),
.A2(n_255),
.B(n_282),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_256),
.B(n_142),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_362),
.B(n_238),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_252),
.B(n_218),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_171),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_228),
.B(n_173),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_369),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_335),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_370),
.Y(n_438)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

BUFx4f_ASAP7_75t_SL g376 ( 
.A(n_369),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_376),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_317),
.A2(n_253),
.B1(n_244),
.B2(n_287),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_377),
.A2(n_388),
.B1(n_389),
.B2(n_358),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_313),
.A2(n_244),
.B1(n_262),
.B2(n_298),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_379),
.A2(n_387),
.B1(n_397),
.B2(n_399),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_381),
.A2(n_410),
.B(n_416),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_309),
.B(n_290),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_398),
.Y(n_426)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_384),
.Y(n_420)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_313),
.A2(n_317),
.B1(n_359),
.B2(n_363),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_317),
.A2(n_173),
.B1(n_262),
.B2(n_204),
.Y(n_388)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_390),
.Y(n_422)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

BUFx24_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_393),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_257),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_394),
.B(n_396),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_349),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_395),
.B(n_406),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_257),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_327),
.A2(n_239),
.B1(n_259),
.B2(n_231),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_310),
.B(n_300),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_327),
.A2(n_353),
.B1(n_326),
.B2(n_345),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_340),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_296),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_405),
.Y(n_443)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_239),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_238),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_312),
.B(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_409),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_332),
.B(n_234),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_413),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_346),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_418),
.Y(n_447)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

A2O1A1Ixp33_ASAP7_75t_SL g428 ( 
.A1(n_415),
.A2(n_351),
.B(n_356),
.C(n_229),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_313),
.A2(n_204),
.B1(n_212),
.B2(n_193),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_335),
.B1(n_336),
.B2(n_333),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_421),
.A2(n_430),
.B1(n_441),
.B2(n_445),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_SL g470 ( 
.A1(n_428),
.A2(n_376),
.B(n_411),
.C(n_416),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_334),
.B1(n_326),
.B2(n_320),
.Y(n_430)
);

OAI22x1_ASAP7_75t_L g431 ( 
.A1(n_379),
.A2(n_315),
.B1(n_354),
.B2(n_322),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_431),
.A2(n_416),
.B1(n_410),
.B2(n_393),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_383),
.A2(n_354),
.B(n_316),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_437),
.A2(n_458),
.B(n_378),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_396),
.A2(n_354),
.B1(n_328),
.B2(n_364),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_371),
.B(n_347),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_450),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_371),
.B(n_338),
.Y(n_450)
);

AOI32xp33_ASAP7_75t_L g451 ( 
.A1(n_380),
.A2(n_360),
.A3(n_352),
.B1(n_368),
.B2(n_338),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_386),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_381),
.A2(n_325),
.B(n_366),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_453),
.A2(n_390),
.B(n_293),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_367),
.C(n_366),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_459),
.C(n_409),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_376),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_380),
.B(n_342),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_398),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_396),
.A2(n_367),
.B(n_325),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_311),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_447),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_462),
.Y(n_515)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_463),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_421),
.A2(n_386),
.B1(n_394),
.B2(n_377),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_464),
.A2(n_442),
.B1(n_435),
.B2(n_438),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_465),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_419),
.B(n_402),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_466),
.B(n_476),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_467),
.B(n_475),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_430),
.A2(n_388),
.B1(n_386),
.B2(n_394),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_468),
.A2(n_479),
.B1(n_433),
.B2(n_453),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_480),
.Y(n_499)
);

AO21x2_ASAP7_75t_SL g521 ( 
.A1(n_470),
.A2(n_428),
.B(n_422),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_471),
.A2(n_495),
.B(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_405),
.Y(n_472)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_410),
.C(n_393),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_486),
.C(n_455),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_404),
.Y(n_474)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_419),
.B(n_357),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_427),
.Y(n_477)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_457),
.Y(n_478)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_429),
.A2(n_417),
.B1(n_370),
.B2(n_408),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_357),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_423),
.B(n_346),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_489),
.Y(n_512)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_447),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_483),
.B(n_488),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_SL g484 ( 
.A(n_436),
.B(n_411),
.C(n_384),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_441),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_444),
.B(n_370),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_493),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_392),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_344),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_344),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_494),
.Y(n_523)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

XOR2x1_ASAP7_75t_L g492 ( 
.A(n_426),
.B(n_384),
.Y(n_492)
);

NOR4xp25_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_428),
.C(n_434),
.D(n_425),
.Y(n_527)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_422),
.B(n_432),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_449),
.A2(n_385),
.B1(n_375),
.B2(n_384),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_414),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_497),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_501),
.A2(n_505),
.B1(n_509),
.B2(n_528),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_461),
.A2(n_446),
.B1(n_436),
.B2(n_420),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_461),
.A2(n_446),
.B1(n_420),
.B2(n_431),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_491),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_511),
.A2(n_521),
.B(n_527),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_485),
.B(n_460),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_472),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_474),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_525),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_462),
.A2(n_438),
.B1(n_435),
.B2(n_442),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_519),
.A2(n_524),
.B1(n_526),
.B2(n_482),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_467),
.B(n_439),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_440),
.B1(n_439),
.B2(n_452),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_468),
.A2(n_440),
.B1(n_452),
.B2(n_434),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_460),
.B(n_425),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_529),
.B(n_531),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_497),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_497),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_534),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_486),
.B(n_361),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_504),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_535),
.B(n_541),
.Y(n_578)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_511),
.A2(n_471),
.B1(n_478),
.B2(n_479),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_537),
.A2(n_548),
.B1(n_521),
.B2(n_508),
.Y(n_574)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_522),
.Y(n_539)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_540),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_499),
.A2(n_463),
.B1(n_495),
.B2(n_496),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_543),
.A2(n_556),
.B1(n_521),
.B2(n_524),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_475),
.C(n_465),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_545),
.C(n_554),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_520),
.B(n_473),
.C(n_484),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_492),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_547),
.B(n_549),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_511),
.A2(n_464),
.B1(n_488),
.B2(n_470),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_505),
.B(n_493),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_558),
.Y(n_582)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_522),
.Y(n_553)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_487),
.C(n_456),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_507),
.B(n_503),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_555),
.B(n_532),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_501),
.A2(n_470),
.B1(n_456),
.B2(n_428),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_516),
.B(n_414),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_557),
.B(n_560),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_513),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_513),
.B(n_470),
.C(n_283),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_564),
.C(n_565),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_507),
.B(n_372),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_532),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_561),
.B(n_503),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_470),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_562),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_500),
.B(n_428),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_521),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_514),
.B(n_264),
.C(n_342),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_514),
.B(n_301),
.C(n_415),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_527),
.A2(n_318),
.B(n_272),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_567),
.A2(n_521),
.B(n_526),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_569),
.A2(n_575),
.B1(n_556),
.B2(n_535),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_585),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_574),
.A2(n_581),
.B1(n_583),
.B2(n_594),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_550),
.A2(n_517),
.B1(n_500),
.B2(n_502),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_506),
.C(n_531),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_576),
.B(n_584),
.Y(n_599)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_537),
.A2(n_508),
.B1(n_498),
.B2(n_502),
.Y(n_581)
);

OAI21xp33_ASAP7_75t_L g584 ( 
.A1(n_545),
.A2(n_523),
.B(n_533),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_498),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_546),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_586),
.B(n_588),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_547),
.B(n_506),
.C(n_528),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_515),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_589),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_542),
.B(n_519),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_552),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_585),
.B(n_554),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_595),
.B(n_605),
.Y(n_628)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_596),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_583),
.A2(n_566),
.B(n_562),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_597),
.A2(n_572),
.B(n_581),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_590),
.A2(n_558),
.B1(n_548),
.B2(n_550),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_598),
.A2(n_606),
.B1(n_608),
.B2(n_574),
.Y(n_617)
);

INVx13_ASAP7_75t_L g603 ( 
.A(n_575),
.Y(n_603)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_603),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_570),
.B(n_549),
.C(n_565),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_604),
.B(n_607),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_590),
.A2(n_536),
.B1(n_559),
.B2(n_566),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_570),
.B(n_564),
.C(n_563),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_593),
.A2(n_567),
.B1(n_518),
.B2(n_297),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_518),
.C(n_260),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_611),
.C(n_616),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_267),
.C(n_226),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_578),
.Y(n_612)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_612),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_578),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_568),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_573),
.B(n_592),
.Y(n_615)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_615),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_276),
.C(n_275),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_617),
.B(n_624),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_614),
.B(n_609),
.Y(n_618)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_618),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_615),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_620),
.Y(n_639)
);

CKINVDCx14_ASAP7_75t_R g620 ( 
.A(n_599),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_602),
.B(n_582),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_598),
.B(n_605),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_626),
.B(n_627),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_604),
.B(n_571),
.C(n_577),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_571),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_185),
.Y(n_650)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_612),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_633),
.B(n_634),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_587),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_597),
.A2(n_568),
.B(n_577),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_635),
.A2(n_601),
.B(n_600),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_637),
.B(n_643),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_632),
.A2(n_596),
.B1(n_606),
.B2(n_608),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_640),
.B(n_642),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_607),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_641),
.B(n_648),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_630),
.B(n_602),
.C(n_610),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_623),
.A2(n_603),
.B1(n_591),
.B2(n_579),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_644),
.B(n_645),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_627),
.B(n_611),
.C(n_616),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_621),
.B(n_591),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_622),
.A2(n_579),
.B(n_193),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_649),
.A2(n_271),
.B(n_242),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_650),
.B(n_651),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_628),
.B(n_185),
.C(n_183),
.Y(n_651)
);

NOR4xp25_ASAP7_75t_L g652 ( 
.A(n_647),
.B(n_618),
.C(n_639),
.D(n_638),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_SL g667 ( 
.A1(n_652),
.A2(n_229),
.B(n_272),
.C(n_232),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_623),
.C(n_631),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_655),
.B(n_659),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_637),
.A2(n_631),
.B1(n_629),
.B2(n_633),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_660),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_648),
.B(n_628),
.C(n_624),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_646),
.A2(n_625),
.B1(n_635),
.B2(n_233),
.Y(n_660)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_662),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_636),
.B(n_286),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_663),
.B(n_281),
.Y(n_668)
);

AOI322xp5_ASAP7_75t_L g664 ( 
.A1(n_653),
.A2(n_643),
.A3(n_644),
.B1(n_636),
.B2(n_642),
.C1(n_645),
.C2(n_650),
.Y(n_664)
);

AO21x1_ASAP7_75t_L g674 ( 
.A1(n_664),
.A2(n_656),
.B(n_654),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_657),
.B(n_651),
.Y(n_666)
);

AOI21xp33_ASAP7_75t_L g676 ( 
.A1(n_666),
.A2(n_661),
.B(n_655),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_SL g672 ( 
.A1(n_667),
.A2(n_229),
.B(n_232),
.C(n_656),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_668),
.B(n_671),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g671 ( 
.A(n_659),
.B(n_183),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_672),
.B(n_674),
.Y(n_679)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_670),
.B(n_654),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_673),
.B(n_676),
.C(n_18),
.Y(n_678)
);

AOI322xp5_ASAP7_75t_L g677 ( 
.A1(n_675),
.A2(n_666),
.A3(n_665),
.B1(n_669),
.B2(n_16),
.C1(n_18),
.C2(n_15),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_677),
.B(n_678),
.C(n_679),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_680),
.B(n_13),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_681),
.B(n_15),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_SL g683 ( 
.A(n_682),
.B(n_15),
.C(n_16),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_683),
.A2(n_16),
.B(n_0),
.Y(n_684)
);


endmodule