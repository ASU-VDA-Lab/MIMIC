module real_aes_7808_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_0), .A2(n_221), .B(n_225), .C(n_262), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_1), .A2(n_216), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_2), .B(n_239), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g199 ( .A(n_4), .Y(n_199) );
AND2x6_ASAP7_75t_L g221 ( .A(n_4), .B(n_197), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_4), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g249 ( .A(n_5), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_6), .A2(n_73), .B1(n_169), .B2(n_173), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_7), .B(n_230), .Y(n_266) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_24), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g214 ( .A(n_9), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_10), .A2(n_250), .B(n_275), .C(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_11), .B(n_239), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_12), .A2(n_53), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_12), .Y(n_183) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_13), .A2(n_26), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_14), .B(n_335), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_15), .A2(n_229), .B(n_231), .C(n_235), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_16), .B(n_230), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_17), .B(n_230), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g295 ( .A(n_18), .Y(n_295) );
INVx1_ASAP7_75t_L g309 ( .A(n_19), .Y(n_309) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_20), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_21), .Y(n_259) );
INVx1_ASAP7_75t_L g332 ( .A(n_22), .Y(n_332) );
INVx2_ASAP7_75t_L g219 ( .A(n_23), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_25), .Y(n_269) );
OAI221xp5_ASAP7_75t_L g190 ( .A1(n_26), .A2(n_41), .B1(n_52), .B2(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g193 ( .A(n_26), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_27), .A2(n_229), .B(n_288), .C(n_290), .Y(n_287) );
INVxp67_ASAP7_75t_L g333 ( .A(n_28), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_29), .A2(n_80), .B1(n_176), .B2(n_177), .Y(n_79) );
INVx1_ASAP7_75t_L g176 ( .A(n_29), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_29), .A2(n_225), .B(n_308), .C(n_314), .Y(n_307) );
CKINVDCx14_ASAP7_75t_R g286 ( .A(n_30), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_30), .A2(n_80), .B1(n_177), .B2(n_286), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_31), .A2(n_80), .B1(n_177), .B2(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_31), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_32), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_33), .A2(n_247), .B(n_248), .C(n_251), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_34), .A2(n_62), .B1(n_141), .B2(n_145), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_35), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_36), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_37), .A2(n_54), .B1(n_161), .B2(n_165), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_38), .A2(n_179), .B1(n_180), .B2(n_186), .Y(n_178) );
INVx1_ASAP7_75t_L g186 ( .A(n_38), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_39), .Y(n_119) );
INVx1_ASAP7_75t_L g223 ( .A(n_40), .Y(n_223) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_41), .A2(n_65), .B1(n_90), .B2(n_94), .Y(n_99) );
INVxp67_ASAP7_75t_L g194 ( .A(n_41), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_42), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_43), .Y(n_100) );
INVx1_ASAP7_75t_L g197 ( .A(n_44), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_45), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_46), .Y(n_126) );
INVx1_ASAP7_75t_L g213 ( .A(n_47), .Y(n_213) );
INVx1_ASAP7_75t_SL g289 ( .A(n_48), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_49), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_50), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g298 ( .A(n_51), .Y(n_298) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_52), .A2(n_69), .B1(n_90), .B2(n_91), .Y(n_97) );
INVx1_ASAP7_75t_L g184 ( .A(n_53), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_55), .A2(n_216), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_56), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_57), .A2(n_216), .B(n_272), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_58), .A2(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g273 ( .A(n_59), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_60), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_61), .A2(n_181), .B1(n_182), .B2(n_185), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_61), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_63), .A2(n_216), .B(n_222), .Y(n_215) );
INVx1_ASAP7_75t_L g276 ( .A(n_64), .Y(n_276) );
INVx2_ASAP7_75t_L g211 ( .A(n_66), .Y(n_211) );
INVx1_ASAP7_75t_L g263 ( .A(n_67), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_68), .A2(n_225), .B(n_297), .C(n_300), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_70), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_71), .B(n_209), .Y(n_253) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
INVx2_ASAP7_75t_L g232 ( .A(n_74), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_75), .A2(n_76), .B1(n_149), .B2(n_154), .Y(n_148) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_187), .B1(n_200), .B2(n_506), .C(n_509), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_178), .Y(n_78) );
INVx1_ASAP7_75t_L g177 ( .A(n_80), .Y(n_177) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_138), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_104), .C(n_125), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_100), .B2(n_101), .Y(n_82) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
INVx2_ASAP7_75t_L g164 ( .A(n_87), .Y(n_164) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g103 ( .A(n_88), .B(n_93), .Y(n_103) );
AND2x2_ASAP7_75t_L g144 ( .A(n_88), .B(n_110), .Y(n_144) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g111 ( .A(n_89), .B(n_99), .Y(n_111) );
AND2x2_ASAP7_75t_L g116 ( .A(n_89), .B(n_93), .Y(n_116) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx2_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
INVx1_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_96), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g147 ( .A(n_96), .B(n_144), .Y(n_147) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g109 ( .A(n_97), .Y(n_109) );
INVx1_ASAP7_75t_L g118 ( .A(n_97), .Y(n_118) );
INVx1_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_97), .B(n_99), .Y(n_158) );
AND2x2_ASAP7_75t_L g117 ( .A(n_98), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g153 ( .A(n_99), .B(n_137), .Y(n_153) );
BUFx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g152 ( .A(n_103), .B(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g167 ( .A(n_103), .B(n_117), .Y(n_167) );
OAI222xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_112), .B1(n_113), .B2(n_119), .C1(n_120), .C2(n_124), .Y(n_104) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
INVx1_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
AND2x4_ASAP7_75t_L g122 ( .A(n_111), .B(n_123), .Y(n_122) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_111), .B(n_129), .Y(n_128) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx1_ASAP7_75t_L g134 ( .A(n_116), .Y(n_134) );
AND2x2_ASAP7_75t_L g143 ( .A(n_117), .B(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g163 ( .A(n_117), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_159), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_148), .Y(n_139) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g172 ( .A(n_144), .B(n_153), .Y(n_172) );
AND2x4_ASAP7_75t_L g174 ( .A(n_144), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx4f_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx6_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
OR2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx1_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_160), .B(n_168), .Y(n_159) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
INVx11_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx6_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_182), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
AND3x1_ASAP7_75t_SL g189 ( .A(n_190), .B(n_195), .C(n_198), .Y(n_189) );
INVxp67_ASAP7_75t_L g514 ( .A(n_190), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
INVx1_ASAP7_75t_SL g515 ( .A(n_195), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_195), .A2(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g526 ( .A(n_195), .Y(n_526) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_196), .B(n_199), .Y(n_520) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_198), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_432), .Y(n_202) );
NOR4xp25_ASAP7_75t_L g203 ( .A(n_204), .B(n_374), .C(n_404), .D(n_414), .Y(n_203) );
OAI211xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_279), .B(n_337), .C(n_364), .Y(n_204) );
OAI222xp33_ASAP7_75t_L g459 ( .A1(n_205), .A2(n_379), .B1(n_460), .B2(n_461), .C1(n_462), .C2(n_463), .Y(n_459) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_254), .Y(n_205) );
AOI33xp33_ASAP7_75t_L g385 ( .A1(n_206), .A2(n_372), .A3(n_373), .B1(n_386), .B2(n_391), .B3(n_393), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_206), .A2(n_443), .B(n_445), .C(n_447), .Y(n_442) );
OR2x2_ASAP7_75t_L g458 ( .A(n_206), .B(n_444), .Y(n_458) );
INVx1_ASAP7_75t_L g491 ( .A(n_206), .Y(n_491) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_241), .Y(n_206) );
INVx2_ASAP7_75t_L g368 ( .A(n_207), .Y(n_368) );
AND2x2_ASAP7_75t_L g384 ( .A(n_207), .B(n_270), .Y(n_384) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_207), .Y(n_419) );
AND2x2_ASAP7_75t_L g448 ( .A(n_207), .B(n_241), .Y(n_448) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_215), .B(n_238), .Y(n_207) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_208), .A2(n_271), .B(n_278), .Y(n_270) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_208), .A2(n_284), .B(n_292), .Y(n_283) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx4_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g325 ( .A(n_210), .Y(n_325) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_211), .B(n_212), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
BUFx2_ASAP7_75t_L g327 ( .A(n_216), .Y(n_327) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_217), .B(n_221), .Y(n_260) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g226 ( .A(n_219), .Y(n_226) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
INVx1_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_220), .Y(n_234) );
INVx3_ASAP7_75t_L g250 ( .A(n_220), .Y(n_250) );
INVx4_ASAP7_75t_SL g237 ( .A(n_221), .Y(n_237) );
BUFx3_ASAP7_75t_L g314 ( .A(n_221), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B(n_228), .C(n_237), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_224), .A2(n_237), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_224), .A2(n_237), .B(n_273), .C(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_224), .A2(n_237), .B(n_286), .C(n_287), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_224), .A2(n_237), .B(n_329), .C(n_330), .Y(n_328) );
INVx5_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
BUFx3_ASAP7_75t_L g252 ( .A(n_226), .Y(n_252) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_226), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_229), .B(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g247 ( .A(n_230), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_233), .B(n_276), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_233), .A2(n_310), .B1(n_332), .B2(n_333), .Y(n_331) );
INVx4_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_237), .B(n_312), .Y(n_508) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_240), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_240), .A2(n_294), .B(n_301), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_240), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g348 ( .A(n_241), .Y(n_348) );
BUFx3_ASAP7_75t_L g356 ( .A(n_241), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_241), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g367 ( .A(n_241), .B(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_241), .B(n_255), .Y(n_396) );
AND2x2_ASAP7_75t_L g465 ( .A(n_241), .B(n_399), .Y(n_465) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_253), .Y(n_241) );
INVx1_ASAP7_75t_L g257 ( .A(n_242), .Y(n_257) );
INVx2_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_242), .A2(n_260), .B(n_306), .C(n_307), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx5_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
INVx2_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g277 ( .A(n_252), .Y(n_277) );
INVx2_ASAP7_75t_SL g359 ( .A(n_254), .Y(n_359) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_270), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_255), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
AND2x2_ASAP7_75t_L g412 ( .A(n_255), .B(n_368), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_255), .B(n_397), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_255), .B(n_399), .Y(n_444) );
AND2x2_ASAP7_75t_L g503 ( .A(n_255), .B(n_448), .Y(n_503) );
INVx4_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g373 ( .A(n_256), .B(n_270), .Y(n_373) );
AND2x2_ASAP7_75t_L g383 ( .A(n_256), .B(n_384), .Y(n_383) );
BUFx3_ASAP7_75t_L g405 ( .A(n_256), .Y(n_405) );
AND3x2_ASAP7_75t_L g464 ( .A(n_256), .B(n_465), .C(n_466), .Y(n_464) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_268), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_261), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_260), .A2(n_295), .B(n_296), .Y(n_294) );
O2A1O1Ixp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_266), .C(n_267), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_264), .A2(n_267), .B(n_298), .C(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_264), .Y(n_507) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_270), .Y(n_355) );
INVx1_ASAP7_75t_SL g399 ( .A(n_270), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_270), .B(n_348), .C(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_317), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_280), .A2(n_383), .B(n_435), .C(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_304), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_282), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_SL g451 ( .A(n_282), .Y(n_451) );
AND2x2_ASAP7_75t_L g472 ( .A(n_282), .B(n_319), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_282), .B(n_381), .Y(n_500) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_293), .Y(n_282) );
AND2x2_ASAP7_75t_L g345 ( .A(n_283), .B(n_336), .Y(n_345) );
INVx2_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
AND2x2_ASAP7_75t_L g372 ( .A(n_283), .B(n_319), .Y(n_372) );
AND2x2_ASAP7_75t_L g422 ( .A(n_283), .B(n_304), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_283), .Y(n_426) );
OAI322xp33_ASAP7_75t_L g509 ( .A1(n_289), .A2(n_510), .A3(n_511), .B1(n_515), .B2(n_516), .C1(n_521), .C2(n_523), .Y(n_509) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g336 ( .A(n_293), .Y(n_336) );
BUFx2_ASAP7_75t_L g362 ( .A(n_293), .Y(n_362) );
AND2x2_ASAP7_75t_L g489 ( .A(n_293), .B(n_304), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
INVx3_ASAP7_75t_SL g319 ( .A(n_304), .Y(n_319) );
AND2x2_ASAP7_75t_L g344 ( .A(n_304), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g351 ( .A(n_304), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g381 ( .A(n_304), .B(n_341), .Y(n_381) );
OR2x2_ASAP7_75t_L g390 ( .A(n_304), .B(n_336), .Y(n_390) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_304), .Y(n_408) );
AND2x2_ASAP7_75t_L g413 ( .A(n_304), .B(n_366), .Y(n_413) );
AND2x2_ASAP7_75t_L g441 ( .A(n_304), .B(n_321), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_304), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g479 ( .A(n_304), .B(n_320), .Y(n_479) );
OR2x6_ASAP7_75t_L g304 ( .A(n_305), .B(n_315), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B(n_311), .C(n_312), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_312), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_313), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g403 ( .A(n_319), .B(n_352), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_319), .B(n_345), .Y(n_431) );
AND2x2_ASAP7_75t_L g449 ( .A(n_319), .B(n_366), .Y(n_449) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_336), .Y(n_320) );
AND2x2_ASAP7_75t_L g350 ( .A(n_321), .B(n_336), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_321), .B(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g388 ( .A(n_321), .Y(n_388) );
OR2x2_ASAP7_75t_L g436 ( .A(n_321), .B(n_356), .Y(n_436) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_326), .B(n_334), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_323), .A2(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g342 ( .A(n_326), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_334), .Y(n_343) );
AND2x2_ASAP7_75t_L g371 ( .A(n_336), .B(n_341), .Y(n_371) );
INVx1_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
AND2x2_ASAP7_75t_L g474 ( .A(n_336), .B(n_352), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_346), .B1(n_349), .B2(n_353), .C1(n_357), .C2(n_360), .Y(n_337) );
INVx1_ASAP7_75t_L g469 ( .A(n_338), .Y(n_469) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_344), .Y(n_338) );
AND2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_345), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_339), .B(n_367), .Y(n_392) );
OAI222xp33_ASAP7_75t_L g414 ( .A1(n_339), .A2(n_415), .B1(n_420), .B2(n_421), .C1(n_429), .C2(n_431), .Y(n_414) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g402 ( .A(n_341), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_341), .B(n_422), .Y(n_462) );
AND2x2_ASAP7_75t_L g473 ( .A(n_341), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g481 ( .A(n_344), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_346), .B(n_397), .Y(n_460) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_348), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g418 ( .A(n_348), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx3_ASAP7_75t_L g363 ( .A(n_351), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_351), .A2(n_454), .B(n_457), .C(n_459), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_351), .B(n_388), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_351), .B(n_371), .Y(n_493) );
AND2x2_ASAP7_75t_L g366 ( .A(n_352), .B(n_362), .Y(n_366) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_356), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g445 ( .A(n_356), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g484 ( .A(n_356), .B(n_384), .Y(n_484) );
INVx1_ASAP7_75t_L g496 ( .A(n_356), .Y(n_496) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_359), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g477 ( .A(n_362), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_367), .B(n_369), .C(n_373), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_395), .B1(n_410), .B2(n_413), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_366), .B(n_380), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_366), .B(n_388), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_367), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g430 ( .A(n_367), .Y(n_430) );
AND2x2_ASAP7_75t_L g437 ( .A(n_367), .B(n_417), .Y(n_437) );
INVx2_ASAP7_75t_L g398 ( .A(n_368), .Y(n_398) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_372), .B(n_376), .C(n_377), .D(n_380), .Y(n_375) );
INVx1_ASAP7_75t_SL g446 ( .A(n_373), .Y(n_446) );
AND2x2_ASAP7_75t_L g490 ( .A(n_373), .B(n_491), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_382), .B(n_385), .C(n_394), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_381), .B(n_451), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_383), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
INVx1_ASAP7_75t_SL g456 ( .A(n_384), .Y(n_456) );
AND2x2_ASAP7_75t_L g495 ( .A(n_384), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_388), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_392), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_393), .B(n_418), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_400), .B(n_402), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g470 ( .A(n_397), .Y(n_470) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx2_ASAP7_75t_L g498 ( .A(n_398), .Y(n_498) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_399), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_409), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_405), .Y(n_417) );
OR2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_SL g450 ( .A1(n_408), .A2(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_439), .B1(n_442), .B2(n_449), .C(n_450), .Y(n_438) );
INVx1_ASAP7_75t_SL g482 ( .A(n_413), .Y(n_482) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g429 ( .A(n_417), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g466 ( .A(n_419), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_426), .B2(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_425), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR4xp25_ASAP7_75t_L g432 ( .A(n_433), .B(n_467), .C(n_480), .D(n_492), .Y(n_432) );
NAND3xp33_ASAP7_75t_SL g433 ( .A(n_434), .B(n_438), .C(n_453), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_436), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_443), .B(n_448), .Y(n_452) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI221xp5_ASAP7_75t_SL g480 ( .A1(n_455), .A2(n_481), .B1(n_482), .B2(n_483), .C(n_485), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_457), .A2(n_472), .B(n_473), .C(n_475), .Y(n_471) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_458), .A2(n_476), .B1(n_478), .B2(n_479), .Y(n_475) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_470), .C(n_471), .Y(n_467) );
INVx1_ASAP7_75t_L g486 ( .A(n_479), .Y(n_486) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_487), .B(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI221xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_494), .B1(n_497), .B2(n_499), .C(n_501), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g519 ( .A(n_507), .Y(n_519) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
endmodule