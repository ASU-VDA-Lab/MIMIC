module fake_aes_280_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
AO31x2_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_5) );
O2A1O1Ixp33_ASAP7_75t_SL g6 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_5), .B(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_8), .B(n_5), .Y(n_9) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .B1(n_6), .B2(n_5), .C(n_2), .Y(n_10) );
NOR3xp33_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .C(n_1), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
NAND5xp2_ASAP7_75t_L g13 ( .A(n_10), .B(n_0), .C(n_1), .D(n_2), .E(n_11), .Y(n_13) );
OA22x2_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_0), .B1(n_2), .B2(n_13), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_12), .Y(n_15) );
endmodule