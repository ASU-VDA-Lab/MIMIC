module fake_jpeg_7965_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_41),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_51),
.B1(n_55),
.B2(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_18),
.B1(n_30),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_53),
.B1(n_58),
.B2(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_30),
.B1(n_18),
.B2(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_32),
.B1(n_33),
.B2(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_20),
.B1(n_17),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_31),
.B1(n_20),
.B2(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_22),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_29),
.B(n_15),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_16),
.C(n_15),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_69),
.B(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_78),
.B(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_85),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_85),
.C(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_47),
.B1(n_50),
.B2(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_22),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_74),
.B1(n_82),
.B2(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_97),
.B1(n_110),
.B2(n_78),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_66),
.B1(n_48),
.B2(n_49),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_97),
.B(n_105),
.C(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_47),
.B1(n_58),
.B2(n_56),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_15),
.Y(n_132)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_73),
.B1(n_35),
.B2(n_15),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_46),
.B(n_57),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_69),
.B(n_106),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_24),
.Y(n_128)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_48),
.B1(n_52),
.B2(n_64),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_118),
.B(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_119),
.B(n_107),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_75),
.B(n_70),
.C(n_72),
.D(n_16),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_70),
.B1(n_80),
.B2(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_127),
.B1(n_130),
.B2(n_104),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_15),
.B(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_93),
.B1(n_89),
.B2(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_93),
.B1(n_107),
.B2(n_102),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_99),
.C(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_142),
.B(n_154),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_155),
.C(n_127),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_115),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_104),
.B(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_88),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_73),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_90),
.B1(n_96),
.B2(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_118),
.B1(n_133),
.B2(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_96),
.B1(n_95),
.B2(n_10),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_156),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_25),
.B1(n_22),
.B2(n_73),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_22),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_130),
.B(n_111),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_166),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_148),
.C(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_139),
.B1(n_133),
.B2(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_124),
.C(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_10),
.C(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_175),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_123),
.Y(n_175)
);

NOR2x1_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_8),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_142),
.B(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_156),
.B1(n_141),
.B2(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_181),
.B1(n_160),
.B2(n_176),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_140),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_183),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_185),
.B(n_176),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_138),
.B1(n_135),
.B2(n_147),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_7),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_112),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_177),
.B1(n_163),
.B2(n_161),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_7),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_9),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_2),
.C(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_194),
.B1(n_178),
.B2(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_210),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_180),
.B(n_157),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_183),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_189),
.C(n_157),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_222),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_210),
.B(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_195),
.C(n_172),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_171),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_198),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_209),
.B(n_200),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_231),
.B1(n_197),
.B2(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_230),
.C(n_220),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_238),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_222),
.C(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_226),
.C(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_207),
.A3(n_202),
.B1(n_6),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_202),
.B1(n_228),
.B2(n_210),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_243),
.A2(n_233),
.B(n_232),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_242),
.A3(n_247),
.B1(n_6),
.B2(n_14),
.C1(n_5),
.C2(n_2),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_246),
.C(n_6),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_14),
.Y(n_252)
);


endmodule