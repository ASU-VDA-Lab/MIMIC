module fake_jpeg_50_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_483;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_60),
.Y(n_198)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_62),
.Y(n_217)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g183 ( 
.A(n_66),
.Y(n_183)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_68),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_75),
.Y(n_139)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_70),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_31),
.B(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_89),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_28),
.B(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_98),
.Y(n_133)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_109),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

BUFx4f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_29),
.B(n_0),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_45),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_125),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

BUFx4f_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

BUFx16f_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_17),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_17),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_54),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_33),
.B(n_0),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_131),
.Y(n_201)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_55),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_138),
.B(n_143),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_140),
.A2(n_194),
.B1(n_41),
.B2(n_30),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_64),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_68),
.A2(n_32),
.B1(n_57),
.B2(n_56),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_146),
.A2(n_150),
.B1(n_20),
.B2(n_50),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_147),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_95),
.A2(n_32),
.B1(n_57),
.B2(n_56),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_65),
.A2(n_58),
.B1(n_52),
.B2(n_49),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_158),
.A2(n_191),
.B1(n_36),
.B2(n_30),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_52),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_161),
.B(n_167),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_40),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_169),
.B(n_172),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_86),
.B(n_40),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_70),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_182),
.B(n_186),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_96),
.B(n_90),
.C(n_80),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_190),
.B(n_114),
.C(n_107),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_76),
.A2(n_33),
.B1(n_38),
.B2(n_49),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_78),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_112),
.B(n_20),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_195),
.B(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_110),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_112),
.B(n_53),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_207),
.B(n_50),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_71),
.B(n_38),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_83),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_221),
.Y(n_254)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_91),
.Y(n_214)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_105),
.B(n_53),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_227),
.Y(n_243)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g222 ( 
.A(n_87),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_71),
.B(n_53),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_107),
.Y(n_260)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_77),
.Y(n_229)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_232),
.Y(n_375)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_233),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g376 ( 
.A(n_234),
.B(n_239),
.C(n_261),
.Y(n_376)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_237),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_244),
.A2(n_263),
.B1(n_268),
.B2(n_269),
.Y(n_337)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_247),
.B(n_293),
.Y(n_366)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_248),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_249),
.A2(n_310),
.B1(n_135),
.B2(n_198),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_164),
.B(n_50),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_255),
.B(n_258),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_256),
.Y(n_368)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_183),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_260),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_134),
.B(n_36),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_262),
.B(n_280),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_166),
.A2(n_94),
.B1(n_92),
.B2(n_77),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_183),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_266),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_267),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_166),
.A2(n_94),
.B1(n_92),
.B2(n_41),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_202),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_168),
.Y(n_270)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_275),
.B1(n_277),
.B2(n_294),
.Y(n_316)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_158),
.A2(n_30),
.B1(n_20),
.B2(n_25),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_201),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_162),
.Y(n_278)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_133),
.B(n_0),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_170),
.Y(n_281)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_1),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_282),
.B(n_284),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_207),
.Y(n_284)
);

OR2x4_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_1),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_285),
.A2(n_150),
.B(n_225),
.Y(n_318)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_208),
.B(n_1),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_287),
.B(n_288),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_149),
.B(n_2),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_160),
.Y(n_289)
);

BUFx4f_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_162),
.Y(n_290)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_292),
.B(n_295),
.Y(n_369)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_188),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_183),
.B(n_3),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_163),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_137),
.B(n_3),
.CI(n_8),
.CON(n_297),
.SN(n_297)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_297),
.B(n_285),
.CI(n_310),
.CON(n_333),
.SN(n_333)
);

AO22x1_ASAP7_75t_SL g298 ( 
.A1(n_144),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_305),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_135),
.B1(n_226),
.B2(n_156),
.Y(n_339)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_176),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_300),
.Y(n_338)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_181),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_301),
.Y(n_350)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_181),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_302),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_319)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_206),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_313),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_141),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_159),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_216),
.A2(n_14),
.B1(n_206),
.B2(n_185),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_216),
.A2(n_185),
.B1(n_223),
.B2(n_199),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_142),
.B(n_177),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_198),
.B(n_175),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_173),
.Y(n_325)
);

OR2x6_ASAP7_75t_SL g423 ( 
.A(n_318),
.B(n_333),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_322),
.A2(n_339),
.B1(n_343),
.B2(n_346),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_349),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_243),
.B(n_177),
.C(n_142),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_364),
.C(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_238),
.B(n_160),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_347),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_271),
.A2(n_157),
.B1(n_193),
.B2(n_153),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_251),
.A2(n_178),
.B1(n_223),
.B2(n_187),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_241),
.B(n_254),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_251),
.A2(n_178),
.A3(n_226),
.B1(n_222),
.B2(n_213),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_250),
.B(n_187),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_354),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_157),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_153),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_357),
.B(n_256),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_247),
.A2(n_224),
.B1(n_145),
.B2(n_165),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_359),
.A2(n_372),
.B1(n_263),
.B2(n_268),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_244),
.A2(n_193),
.B1(n_145),
.B2(n_165),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_367),
.B1(n_371),
.B2(n_246),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_266),
.B(n_171),
.C(n_212),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_294),
.A2(n_224),
.B1(n_171),
.B2(n_212),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_298),
.A2(n_197),
.B1(n_136),
.B2(n_184),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_136),
.B1(n_213),
.B2(n_222),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_252),
.B(n_184),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_308),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

INVx13_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

BUFx2_ASAP7_75t_R g449 ( 
.A(n_383),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_393),
.B1(n_394),
.B2(n_412),
.Y(n_434)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_303),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_386),
.B(n_403),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_361),
.A2(n_278),
.B1(n_290),
.B2(n_245),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_387),
.A2(n_424),
.B(n_248),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_265),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_398),
.Y(n_433)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_389),
.Y(n_438)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_318),
.A2(n_324),
.B(n_337),
.C(n_354),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_391),
.A2(n_377),
.B(n_303),
.Y(n_458)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_324),
.A2(n_269),
.B1(n_232),
.B2(n_281),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_314),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_397),
.B(n_402),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_347),
.B(n_246),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_235),
.C(n_240),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_411),
.C(n_421),
.Y(n_430)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx13_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_410),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_353),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_315),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_405),
.Y(n_429)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_345),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_406),
.B(n_415),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_305),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_408),
.B(n_416),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_357),
.A2(n_237),
.B1(n_301),
.B2(n_274),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_409),
.A2(n_426),
.B1(n_362),
.B2(n_350),
.Y(n_431)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_231),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_322),
.A2(n_272),
.B1(n_253),
.B2(n_291),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_417),
.Y(n_440)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_328),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_328),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_366),
.B(n_293),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_332),
.B(n_259),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_425),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_316),
.A2(n_302),
.B1(n_279),
.B2(n_273),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_331),
.B(n_300),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_363),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_427),
.A2(n_321),
.B1(n_317),
.B2(n_365),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_374),
.B(n_359),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_428),
.A2(n_447),
.B(n_459),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_394),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_402),
.A2(n_333),
.B1(n_342),
.B2(n_319),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_432),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_334),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_437),
.C(n_453),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_364),
.C(n_325),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g443 ( 
.A1(n_414),
.A2(n_333),
.A3(n_358),
.B1(n_349),
.B2(n_372),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_448),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_395),
.A2(n_346),
.B1(n_317),
.B2(n_321),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_446),
.A2(n_464),
.B1(n_467),
.B2(n_393),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_395),
.A2(n_377),
.B(n_336),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_420),
.A2(n_365),
.B1(n_323),
.B2(n_375),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_450),
.A2(n_456),
.B1(n_387),
.B2(n_392),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_452),
.A2(n_368),
.B1(n_307),
.B2(n_283),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_320),
.C(n_330),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_391),
.A2(n_375),
.B1(n_352),
.B2(n_335),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_458),
.A2(n_463),
.B(n_469),
.C(n_344),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_423),
.A2(n_335),
.B(n_360),
.Y(n_459)
);

XOR2x1_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_360),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_414),
.A2(n_270),
.B1(n_257),
.B2(n_242),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_391),
.A2(n_407),
.B1(n_423),
.B2(n_424),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_384),
.A2(n_344),
.B(n_373),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_468),
.Y(n_470)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_468),
.Y(n_472)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_473),
.B(n_475),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_474),
.A2(n_483),
.B1(n_487),
.B2(n_469),
.Y(n_510)
);

OAI32xp33_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_407),
.A3(n_391),
.B1(n_399),
.B2(n_386),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_329),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_476),
.B(n_477),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_373),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_478),
.B(n_505),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_433),
.B(n_421),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_481),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_429),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_486),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_435),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_429),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_467),
.A2(n_412),
.B1(n_427),
.B2(n_404),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_433),
.B(n_419),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_503),
.Y(n_522)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_415),
.Y(n_490)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_490),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_466),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_502),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_436),
.B(n_378),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_441),
.C(n_455),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_413),
.Y(n_493)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_434),
.A2(n_382),
.B1(n_425),
.B2(n_390),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_494),
.A2(n_500),
.B1(n_464),
.B2(n_446),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_437),
.B(n_379),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_497),
.B(n_430),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_498),
.A2(n_459),
.B(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_499),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_434),
.A2(n_406),
.B1(n_400),
.B2(n_385),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_440),
.B(n_444),
.Y(n_501)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_410),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_338),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_381),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_507),
.Y(n_525)
);

INVx13_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_457),
.Y(n_507)
);

INVx13_ASAP7_75t_L g508 ( 
.A(n_449),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_508),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_510),
.A2(n_515),
.B1(n_524),
.B2(n_534),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_473),
.A2(n_432),
.B1(n_431),
.B2(n_450),
.Y(n_515)
);

AO21x1_ASAP7_75t_L g570 ( 
.A1(n_517),
.A2(n_519),
.B(n_498),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_478),
.B(n_458),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_463),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_523),
.B(n_527),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_488),
.A2(n_456),
.B1(n_440),
.B2(n_447),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_457),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_526),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_471),
.B(n_430),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_466),
.B1(n_443),
.B2(n_452),
.Y(n_534)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_536),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_537),
.B(n_494),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_497),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_538),
.B(n_539),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_442),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_540),
.B(n_460),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_490),
.B(n_453),
.Y(n_541)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_470),
.B(n_455),
.Y(n_542)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_542),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_546),
.Y(n_563)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_545),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_495),
.B(n_461),
.Y(n_546)
);

AOI21xp33_ASAP7_75t_L g547 ( 
.A1(n_522),
.A2(n_496),
.B(n_485),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_472),
.Y(n_549)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_549),
.Y(n_580)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_550),
.Y(n_581)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_516),
.Y(n_552)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_553),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_512),
.A2(n_474),
.B1(n_478),
.B2(n_480),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_555),
.A2(n_565),
.B1(n_569),
.B2(n_573),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_513),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_557),
.Y(n_596)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_513),
.A2(n_498),
.B(n_502),
.C(n_491),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_560),
.A2(n_570),
.B(n_531),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_496),
.C(n_495),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_561),
.B(n_564),
.C(n_567),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_486),
.Y(n_562)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_562),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_500),
.C(n_487),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_521),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_499),
.C(n_442),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_489),
.C(n_461),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_571),
.B(n_575),
.C(n_518),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_462),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_572),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_512),
.A2(n_483),
.B1(n_498),
.B2(n_475),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_528),
.B(n_462),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_523),
.B(n_460),
.C(n_505),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_535),
.B(n_498),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_578),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_520),
.A2(n_519),
.B1(n_544),
.B2(n_511),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_577),
.A2(n_579),
.B(n_544),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_519),
.A2(n_466),
.B(n_506),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_558),
.A2(n_531),
.B1(n_517),
.B2(n_514),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_583),
.A2(n_587),
.B1(n_604),
.B2(n_559),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_566),
.B(n_546),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_592),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_586),
.B(n_590),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_577),
.A2(n_532),
.B(n_536),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_569),
.A2(n_511),
.B1(n_514),
.B2(n_532),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_563),
.B(n_525),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_570),
.A2(n_537),
.B(n_545),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_594),
.B(n_599),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_605),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_549),
.B(n_533),
.Y(n_598)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_598),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_573),
.A2(n_533),
.B(n_530),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_567),
.B(n_509),
.C(n_529),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_571),
.C(n_554),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_569),
.A2(n_530),
.B1(n_529),
.B2(n_482),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_SL g605 ( 
.A(n_563),
.B(n_566),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_583),
.A2(n_555),
.B1(n_556),
.B2(n_554),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_606),
.A2(n_609),
.B1(n_617),
.B2(n_624),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_607),
.B(n_610),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_600),
.A2(n_562),
.B1(n_548),
.B2(n_576),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_564),
.C(n_568),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_598),
.Y(n_611)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_611),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_551),
.Y(n_613)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_613),
.Y(n_631)
);

FAx1_ASAP7_75t_SL g614 ( 
.A(n_585),
.B(n_561),
.CI(n_560),
.CON(n_614),
.SN(n_614)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_614),
.B(n_615),
.Y(n_640)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_601),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_616),
.B(n_626),
.Y(n_632)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_581),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_592),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_620),
.B(n_621),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_591),
.B(n_605),
.C(n_568),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_591),
.B(n_575),
.C(n_579),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_622),
.B(n_584),
.C(n_588),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_623),
.A2(n_580),
.B1(n_600),
.B2(n_586),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_552),
.Y(n_624)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_581),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_582),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_582),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_628),
.B(n_642),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_607),
.B(n_603),
.C(n_588),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_630),
.B(n_635),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_612),
.B(n_594),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_644),
.Y(n_648)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_634),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_613),
.B(n_624),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_618),
.A2(n_589),
.B(n_590),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_636),
.A2(n_640),
.B(n_618),
.Y(n_649)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_637),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_610),
.B(n_622),
.C(n_625),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_641),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_625),
.B(n_599),
.C(n_604),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_595),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_595),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_608),
.B(n_550),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_646),
.B(n_627),
.Y(n_647)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_647),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_649),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_643),
.B(n_606),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_655),
.Y(n_672)
);

OAI21x1_ASAP7_75t_SL g654 ( 
.A1(n_631),
.A2(n_626),
.B(n_617),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_654),
.A2(n_637),
.B(n_645),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_639),
.B(n_621),
.C(n_609),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_632),
.A2(n_614),
.B1(n_629),
.B2(n_633),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_659),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_644),
.A2(n_614),
.B1(n_482),
.B2(n_438),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_638),
.B(n_448),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_660),
.B(n_642),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_438),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_661),
.B(n_648),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_664),
.A2(n_665),
.B(n_671),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_656),
.A2(n_651),
.B(n_652),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_666),
.B(n_236),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_SL g667 ( 
.A1(n_658),
.A2(n_630),
.B(n_628),
.C(n_508),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_667),
.A2(n_659),
.B(n_650),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_368),
.C(n_401),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_668),
.B(n_670),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_657),
.A2(n_405),
.B(n_233),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_668),
.B(n_648),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_673),
.B(n_676),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_674),
.A2(n_677),
.B(n_678),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_660),
.C(n_405),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_405),
.Y(n_677)
);

XOR2xp5_ASAP7_75t_L g680 ( 
.A(n_669),
.B(n_383),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_680),
.A2(n_671),
.B(n_389),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_SL g681 ( 
.A1(n_677),
.A2(n_663),
.B(n_667),
.C(n_669),
.Y(n_681)
);

OAI31xp33_ASAP7_75t_SL g685 ( 
.A1(n_681),
.A2(n_682),
.A3(n_675),
.B(n_678),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_685),
.B(n_686),
.C(n_684),
.Y(n_687)
);

AOI322xp5_ASAP7_75t_L g686 ( 
.A1(n_683),
.A2(n_152),
.A3(n_236),
.B1(n_306),
.B2(n_679),
.C1(n_663),
.C2(n_665),
.Y(n_686)
);

AOI21x1_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_236),
.B(n_306),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_688),
.Y(n_689)
);

BUFx24_ASAP7_75t_SL g690 ( 
.A(n_689),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_690),
.B(n_306),
.Y(n_691)
);


endmodule