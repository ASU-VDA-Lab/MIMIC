module real_jpeg_10653_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_0),
.A2(n_11),
.B1(n_13),
.B2(n_17),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_3),
.A2(n_14),
.B1(n_15),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_4),
.A2(n_14),
.B1(n_15),
.B2(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_5),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B1(n_22),
.B2(n_32),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_19),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_11),
.A2(n_13),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);


endmodule