module fake_jpeg_28746_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_52),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_47),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_42),
.B1(n_59),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_74),
.B1(n_47),
.B2(n_41),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_42),
.B1(n_40),
.B2(n_53),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_50),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_63),
.B(n_20),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_80),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_68),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_89),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_45),
.C(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_5),
.C(n_6),
.Y(n_102)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_1),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_79),
.B1(n_77),
.B2(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_104),
.B1(n_19),
.B2(n_21),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_3),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_22),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_11),
.C(n_12),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_107),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_113),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_37),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_101),
.C(n_27),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_101),
.B(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_107),
.B(n_116),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_123),
.B(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_119),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_121),
.B(n_104),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_36),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_26),
.B(n_28),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_35),
.Y(n_132)
);


endmodule