module real_jpeg_12764_n_17 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_3),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_123),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_123),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_123),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_6),
.B(n_30),
.C(n_46),
.Y(n_155)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_6),
.B(n_79),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_114),
.B(n_167),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_6),
.A2(n_60),
.B(n_78),
.C(n_194),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_6),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_6),
.B(n_55),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_41),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_7),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_41),
.B1(n_43),
.B2(n_81),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_81),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_41),
.B1(n_43),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_163),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_163),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_163),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_12),
.A2(n_41),
.B1(n_43),
.B2(n_57),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_41),
.B1(n_43),
.B2(n_70),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_70),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_15),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_15),
.A2(n_40),
.B1(n_55),
.B2(n_56),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_256)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_324),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_311),
.B(n_323),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_139),
.B(n_308),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_126),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_101),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_22),
.B(n_101),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_23),
.B(n_72),
.C(n_87),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_53),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_24),
.A2(n_25),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_26),
.A2(n_27),
.B1(n_53),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_26),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_33),
.B(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_28),
.A2(n_33),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_28),
.B(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_28),
.A2(n_33),
.B1(n_113),
.B2(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_29),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_33),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_35),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_49),
.B2(n_52),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_39),
.A2(n_44),
.B1(n_52),
.B2(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_43),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_41),
.B(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_43),
.A2(n_77),
.B(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_52),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_44),
.B(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_44),
.A2(n_52),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_44),
.A2(n_52),
.B1(n_118),
.B2(n_245),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_50),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_48),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_48),
.B(n_151),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_48),
.A2(n_164),
.B(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_52),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_58),
.B1(n_66),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_63),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_56),
.A2(n_66),
.B(n_151),
.C(n_238),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_56),
.A2(n_60),
.A3(n_63),
.B1(n_239),
.B2(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_66),
.B1(n_99),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_58),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_58),
.A2(n_64),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_58),
.A2(n_66),
.B1(n_122),
.B2(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_59),
.B(n_61),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_65),
.A2(n_219),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_65),
.A2(n_219),
.B1(n_318),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_87),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_73),
.B(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_80),
.B1(n_82),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_82),
.B1(n_92),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_74),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_74),
.A2(n_82),
.B1(n_214),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_74),
.A2(n_200),
.B(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_79),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_75),
.B(n_201),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_75),
.A2(n_79),
.B(n_315),
.Y(n_314)
);

NOR2x1_ASAP7_75t_R g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_79),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_82),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_82),
.A2(n_120),
.B(n_215),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_85),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_85),
.A2(n_152),
.B(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_89),
.B(n_94),
.C(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_94),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_94),
.B(n_131),
.C(n_135),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_98),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_98),
.B(n_130),
.C(n_137),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_107),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_108),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.C(n_121),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_109),
.A2(n_110),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_111),
.A2(n_116),
.B1(n_117),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_111),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_114),
.A2(n_115),
.B1(n_196),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_114),
.A2(n_115),
.B1(n_222),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_115),
.A2(n_173),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_115),
.B(n_151),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_115),
.A2(n_181),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_119),
.B(n_121),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_125),
.B(n_237),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_126),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_127),
.B(n_138),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_132),
.Y(n_317)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_136),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_302),
.B(n_307),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_290),
.B(n_301),
.Y(n_140)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_258),
.A3(n_283),
.B1(n_288),
.B2(n_289),
.C(n_333),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_231),
.B(n_257),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_208),
.B(n_230),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_189),
.B(n_207),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_169),
.B(n_188),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_177),
.B(n_187),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_175),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B(n_186),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_202),
.C(n_206),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_195),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_210),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_223),
.B2(n_224),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_226),
.C(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_217),
.C(n_221),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_247),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_248),
.C(n_249),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_240),
.B2(n_246),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_241),
.C(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_273),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_273),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_269),
.C(n_272),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_261),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_267),
.C(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_272),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_277),
.C(n_282),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_300),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_322),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_322),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_321),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_314),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_319),
.C(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_326),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);


endmodule