module fake_ariane_111_n_604 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_604);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_604;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_22),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_85),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_24),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_50),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_5),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_36),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_20),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_38),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_58),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_21),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_11),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_19),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_66),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_53),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_70),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_69),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_51),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_39),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_16),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_64),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_41),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_62),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_49),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_77),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_90),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_0),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_1),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_151),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_2),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_129),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_131),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_154),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_137),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_142),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_143),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_145),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_138),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_149),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_193),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_171),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_196),
.B(n_157),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_152),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_153),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_192),
.B(n_189),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_197),
.B(n_4),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_234),
.B(n_157),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_200),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_204),
.B(n_155),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_194),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_160),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_161),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_164),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_250),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_166),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_167),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_168),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_253),
.A2(n_173),
.B1(n_185),
.B2(n_179),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_242),
.B(n_170),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_177),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_250),
.B(n_186),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_258),
.A2(n_165),
.B1(n_158),
.B2(n_6),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_158),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_274),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_158),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_256),
.B(n_165),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_165),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_265),
.B(n_4),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_253),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_277),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_277),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_8),
.Y(n_339)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_264),
.B(n_9),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_5),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_268),
.B(n_6),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_267),
.B(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_238),
.B(n_7),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_267),
.B(n_7),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_266),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_313),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_320),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

AND2x6_ASAP7_75t_SL g360 ( 
.A(n_335),
.B(n_280),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

OR2x6_ASAP7_75t_SL g362 ( 
.A(n_337),
.B(n_272),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_262),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_275),
.B1(n_241),
.B2(n_283),
.C(n_266),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_270),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_241),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_282),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_334),
.A2(n_283),
.B1(n_278),
.B2(n_279),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

BUFx6f_ASAP7_75t_SL g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

OAI221xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_275),
.B1(n_270),
.B2(n_273),
.C(n_278),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_277),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_263),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_294),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_302),
.A2(n_276),
.B1(n_282),
.B2(n_281),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_338),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_310),
.B(n_282),
.Y(n_389)
);

AO22x2_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_282),
.B1(n_281),
.B2(n_17),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_281),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_281),
.B1(n_15),
.B2(n_18),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_299),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_127),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_319),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_289),
.B(n_14),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_315),
.B(n_23),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_297),
.B(n_25),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_332),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_350),
.B(n_332),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_369),
.B(n_344),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_388),
.B(n_290),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_311),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_381),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_330),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_330),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_389),
.B(n_298),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_352),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_363),
.B(n_404),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_317),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_404),
.B(n_300),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_333),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_348),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_339),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_399),
.B(n_339),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_377),
.B(n_340),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_339),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_400),
.B(n_339),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_397),
.B(n_27),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_385),
.B(n_29),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_377),
.B(n_30),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_386),
.B(n_402),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_384),
.B(n_31),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_372),
.B(n_32),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_373),
.B(n_33),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_SL g434 ( 
.A(n_405),
.B(n_34),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_35),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_387),
.B(n_37),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_40),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_354),
.B(n_42),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_43),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_45),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_355),
.B(n_46),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_378),
.B(n_358),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_409),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_419),
.A2(n_371),
.B(n_403),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_395),
.B(n_393),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_427),
.B(n_414),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_403),
.B(n_380),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_442),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_375),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_435),
.A2(n_368),
.B(n_396),
.Y(n_450)
);

AO31x2_ASAP7_75t_L g451 ( 
.A1(n_416),
.A2(n_366),
.A3(n_361),
.B(n_364),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_390),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_420),
.A2(n_367),
.B(n_365),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_370),
.B(n_392),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_440),
.A2(n_390),
.B1(n_394),
.B2(n_379),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_407),
.A2(n_360),
.B(n_362),
.C(n_394),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_47),
.B(n_52),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_54),
.B(n_56),
.Y(n_459)
);

OAI22x1_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_410),
.B(n_63),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_67),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_68),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_439),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_433),
.B(n_436),
.Y(n_466)
);

AO32x2_ASAP7_75t_L g467 ( 
.A1(n_408),
.A2(n_126),
.A3(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_443),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_462),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_465),
.Y(n_472)
);

INVx8_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

NOR3xp33_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_406),
.C(n_424),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_468),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_450),
.A2(n_428),
.B(n_425),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_431),
.B(n_429),
.C(n_434),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_426),
.B(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_455),
.B(n_422),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_421),
.Y(n_481)
);

BUFx2_ASAP7_75t_SL g482 ( 
.A(n_448),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_463),
.B(n_422),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_449),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_446),
.A2(n_78),
.B(n_80),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_466),
.A2(n_81),
.B(n_84),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_87),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_125),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_467),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_447),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_459),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_489),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_472),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_472),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_477),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_491),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_473),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_473),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_476),
.A2(n_459),
.B(n_457),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_488),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_474),
.B(n_490),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_490),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_487),
.A2(n_89),
.B(n_91),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_478),
.A2(n_95),
.B(n_99),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_R g521 ( 
.A(n_514),
.B(n_483),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_484),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_483),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_514),
.B(n_100),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_102),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_105),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_R g531 ( 
.A(n_510),
.B(n_107),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_499),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_509),
.B(n_110),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_112),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_506),
.B(n_115),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_116),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_504),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_119),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_509),
.B(n_517),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_517),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_493),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_538),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_526),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_508),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_508),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_533),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_518),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_502),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_501),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_503),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_532),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_540),
.A2(n_494),
.B1(n_520),
.B2(n_493),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_501),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_503),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_512),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_549),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_548),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_555),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_552),
.B(n_524),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_549),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_498),
.Y(n_566)
);

OAI32xp33_ASAP7_75t_L g567 ( 
.A1(n_561),
.A2(n_525),
.A3(n_531),
.B1(n_556),
.B2(n_558),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_565),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_559),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_556),
.C(n_546),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_546),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_566),
.B(n_547),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_562),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_554),
.Y(n_574)
);

CKINVDCx8_ASAP7_75t_R g575 ( 
.A(n_567),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_544),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_569),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_571),
.B(n_545),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_576),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_574),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_578),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_562),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_575),
.B(n_568),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_581),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_579),
.Y(n_585)
);

XNOR2x1_ASAP7_75t_L g586 ( 
.A(n_583),
.B(n_572),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_580),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_585),
.B(n_579),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_587),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_589),
.Y(n_590)
);

AOI221xp5_ASAP7_75t_SL g591 ( 
.A1(n_590),
.A2(n_588),
.B1(n_582),
.B2(n_550),
.C(n_586),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_591),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_592),
.B(n_548),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_593),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_552),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_595),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_596),
.A2(n_534),
.B1(n_535),
.B2(n_516),
.Y(n_597)
);

NAND4xp25_ASAP7_75t_SL g598 ( 
.A(n_597),
.B(n_564),
.C(n_537),
.D(n_529),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_519),
.B(n_529),
.Y(n_599)
);

OAI221xp5_ASAP7_75t_SL g600 ( 
.A1(n_598),
.A2(n_557),
.B1(n_513),
.B2(n_535),
.C(n_521),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_600),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_599),
.Y(n_602)
);

AOI221xp5_ASAP7_75t_L g603 ( 
.A1(n_602),
.A2(n_516),
.B1(n_513),
.B2(n_563),
.C(n_124),
.Y(n_603)
);

AOI211xp5_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_601),
.B(n_516),
.C(n_511),
.Y(n_604)
);


endmodule