module fake_jpeg_2654_n_493 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_49),
.Y(n_155)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_62),
.Y(n_104)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_0),
.Y(n_100)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_60),
.B(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_66),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_67),
.Y(n_156)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_7),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_86),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_94),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_29),
.B1(n_28),
.B2(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_25),
.B1(n_36),
.B2(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_98),
.A2(n_81),
.B1(n_93),
.B2(n_82),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_25),
.B1(n_36),
.B2(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_99),
.A2(n_109),
.B1(n_121),
.B2(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_100),
.B(n_98),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_50),
.A2(n_45),
.B1(n_29),
.B2(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_110),
.B1(n_113),
.B2(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_35),
.B1(n_25),
.B2(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_29),
.B1(n_28),
.B2(n_48),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_29),
.B1(n_28),
.B2(n_48),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_76),
.A2(n_29),
.B1(n_34),
.B2(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_23),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_67),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_139),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_44),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_59),
.A2(n_48),
.B1(n_19),
.B2(n_31),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_149),
.B1(n_152),
.B2(n_77),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_80),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_64),
.B1(n_49),
.B2(n_94),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_52),
.A2(n_43),
.B1(n_41),
.B2(n_34),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_67),
.B1(n_63),
.B2(n_68),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_61),
.A2(n_32),
.B1(n_23),
.B2(n_26),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_84),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_26),
.B1(n_38),
.B2(n_2),
.Y(n_152)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_158),
.Y(n_252)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_163),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_108),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_165),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVxp67_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_54),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_175),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_171),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_153),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_173),
.Y(n_264)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_91),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_176),
.B(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_177),
.B(n_182),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_199),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_56),
.C(n_73),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_185),
.Y(n_240)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_0),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_95),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_64),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_0),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_197),
.Y(n_262)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_193),
.A2(n_196),
.B1(n_198),
.B2(n_209),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_1),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_26),
.B1(n_88),
.B2(n_94),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_111),
.B(n_1),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_154),
.A3(n_147),
.B1(n_103),
.B2(n_122),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_202),
.A2(n_123),
.B(n_124),
.Y(n_219)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_107),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_6),
.Y(n_259)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_103),
.B(n_107),
.C(n_122),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_129),
.C(n_119),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_118),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_1),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_120),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_114),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_214),
.B(n_26),
.C(n_3),
.Y(n_246)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_145),
.B1(n_115),
.B2(n_97),
.Y(n_216)
);

AO21x2_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_223),
.B(n_253),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_219),
.A2(n_174),
.B(n_159),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_97),
.B1(n_142),
.B2(n_102),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_228),
.B1(n_242),
.B2(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_188),
.A2(n_129),
.B1(n_119),
.B2(n_123),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_239),
.B(n_254),
.C(n_173),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_183),
.A2(n_140),
.B1(n_142),
.B2(n_112),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_177),
.A2(n_140),
.B1(n_112),
.B2(n_26),
.Y(n_244)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_175),
.A2(n_26),
.B(n_3),
.C(n_4),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_248),
.A2(n_213),
.B(n_210),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_162),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_249),
.A2(n_256),
.B1(n_182),
.B2(n_195),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_162),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_169),
.B(n_2),
.C(n_6),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_160),
.A2(n_204),
.B1(n_199),
.B2(n_197),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_206),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_172),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_265),
.B(n_269),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_205),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_238),
.A2(n_160),
.B1(n_193),
.B2(n_189),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_273),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_225),
.B(n_256),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_281),
.B(n_289),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_234),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_275),
.B(n_282),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_213),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_202),
.B(n_161),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_234),
.B(n_168),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_290),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_184),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_190),
.B(n_191),
.C(n_192),
.D(n_203),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g345 ( 
.A1(n_288),
.A2(n_309),
.B(n_246),
.C(n_258),
.D(n_230),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_212),
.B(n_200),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_229),
.B(n_211),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_180),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_293),
.Y(n_325)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_157),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_298),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_194),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_301),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_233),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_306),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_214),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_304),
.C(n_240),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_218),
.B(n_9),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_10),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_221),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_307),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_242),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_217),
.B1(n_260),
.B2(n_220),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_13),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_272),
.A2(n_281),
.B1(n_274),
.B2(n_277),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_310),
.A2(n_316),
.B1(n_285),
.B2(n_273),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_263),
.B1(n_228),
.B2(n_227),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_313),
.A2(n_322),
.B1(n_327),
.B2(n_343),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_272),
.A2(n_244),
.B1(n_238),
.B2(n_241),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_306),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_222),
.C(n_257),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_323),
.C(n_344),
.Y(n_357)
);

AOI22x1_ASAP7_75t_SL g322 ( 
.A1(n_285),
.A2(n_248),
.B1(n_246),
.B2(n_257),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_245),
.C(n_231),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_272),
.A2(n_298),
.B1(n_292),
.B2(n_287),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_273),
.A2(n_237),
.B1(n_236),
.B2(n_264),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_272),
.A2(n_249),
.B1(n_217),
.B2(n_247),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_258),
.C(n_237),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_348),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_230),
.C(n_260),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_289),
.C(n_300),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_304),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_282),
.Y(n_351)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_371),
.B(n_379),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_312),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_285),
.B(n_291),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_364),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_355),
.B(n_356),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_266),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_265),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_366),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_317),
.A2(n_285),
.B1(n_268),
.B2(n_293),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_359),
.A2(n_361),
.B1(n_370),
.B2(n_324),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_369),
.C(n_378),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_317),
.A2(n_268),
.B1(n_291),
.B2(n_288),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_310),
.A2(n_308),
.B1(n_267),
.B2(n_279),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_365),
.A2(n_374),
.B1(n_380),
.B2(n_324),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_296),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_325),
.B(n_278),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_319),
.B(n_271),
.C(n_294),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_329),
.A2(n_283),
.B1(n_280),
.B2(n_301),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_329),
.A2(n_246),
.B(n_302),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_299),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_323),
.B(n_220),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_373),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_307),
.B1(n_221),
.B2(n_16),
.Y(n_374)
);

OAI32xp33_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_315),
.A3(n_347),
.B1(n_330),
.B2(n_320),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_377),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_318),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_13),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_315),
.A2(n_13),
.B(n_15),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_313),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_324),
.B(n_326),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_385),
.A2(n_15),
.B(n_16),
.Y(n_429)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_346),
.C(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_401),
.C(n_404),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_389),
.A2(n_391),
.B1(n_348),
.B2(n_379),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_316),
.B1(n_336),
.B2(n_318),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_312),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_375),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_352),
.A2(n_339),
.B1(n_345),
.B2(n_336),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_394),
.A2(n_407),
.B1(n_359),
.B2(n_361),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_376),
.A2(n_321),
.B1(n_322),
.B2(n_340),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_354),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_406),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_351),
.A2(n_333),
.A3(n_342),
.B1(n_340),
.B2(n_314),
.Y(n_398)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_367),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_399),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_321),
.C(n_342),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_331),
.C(n_338),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_331),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_365),
.A2(n_349),
.B1(n_364),
.B2(n_367),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_389),
.A2(n_349),
.B1(n_377),
.B2(n_376),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_414),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_424),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_425),
.B1(n_430),
.B2(n_391),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_403),
.A2(n_380),
.B1(n_374),
.B2(n_371),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_360),
.C(n_372),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_421),
.C(n_423),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_405),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_422),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_429),
.Y(n_447)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_420),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_363),
.C(n_370),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_402),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_378),
.C(n_338),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_356),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_314),
.C(n_333),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_427),
.C(n_406),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_332),
.C(n_362),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_390),
.Y(n_434)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_SL g432 ( 
.A(n_413),
.B(n_403),
.C(n_387),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_435),
.C(n_437),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_381),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_SL g437 ( 
.A(n_430),
.B(n_393),
.C(n_383),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_410),
.B(n_393),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_448),
.Y(n_456)
);

A2O1A1O1Ixp25_ASAP7_75t_L g440 ( 
.A1(n_411),
.A2(n_385),
.B(n_400),
.C(n_392),
.D(n_383),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_440),
.A2(n_382),
.B(n_429),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_414),
.B1(n_386),
.B2(n_382),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_410),
.B(n_384),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_442),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_397),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_444),
.C(n_445),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_407),
.C(n_396),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_426),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_394),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_419),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_460),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_420),
.B1(n_419),
.B2(n_408),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_452),
.A2(n_462),
.B1(n_449),
.B2(n_428),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_433),
.A2(n_417),
.B(n_409),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_455),
.A2(n_457),
.B(n_447),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_433),
.A2(n_417),
.B(n_408),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_431),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_423),
.C(n_412),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_445),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_437),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_432),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_464),
.A2(n_465),
.B(n_467),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_440),
.B(n_447),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_458),
.B(n_444),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_472),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_451),
.B1(n_454),
.B2(n_462),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_439),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_443),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_457),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_466),
.B(n_456),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_480),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_476),
.A2(n_467),
.B(n_461),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_481),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_477),
.A2(n_465),
.B(n_453),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_483),
.B(n_477),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_478),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_487),
.B(n_479),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_486),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_488),
.A2(n_489),
.B1(n_474),
.B2(n_482),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_460),
.Y(n_491)
);

AOI32xp33_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_453),
.A3(n_473),
.B1(n_439),
.B2(n_17),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_17),
.Y(n_493)
);


endmodule