module fake_netlist_5_2223_n_193 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_193);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_193;

wire n_137;
wire n_168;
wire n_164;
wire n_191;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_98;
wire n_66;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_123;
wire n_38;
wire n_139;
wire n_113;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_154;
wire n_62;
wire n_138;
wire n_148;
wire n_100;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_170;
wire n_162;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_115;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVxp33_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_4),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_52),
.B1(n_35),
.B2(n_41),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_53),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_46),
.B1(n_45),
.B2(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_38),
.Y(n_78)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_55),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

OAI221xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_31),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_11),
.B1(n_12),
.B2(n_21),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_22),
.B(n_24),
.C(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_55),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx8_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_64),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_78),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_75),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_75),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_91),
.B(n_86),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_89),
.B(n_93),
.C(n_78),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_89),
.B(n_82),
.C(n_67),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_94),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_95),
.B(n_97),
.Y(n_113)
);

NOR2x1_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_104),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_101),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_102),
.B(n_98),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_79),
.B(n_94),
.Y(n_121)
);

AOI211xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_70),
.B(n_110),
.C(n_72),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_101),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_115),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_127),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_117),
.B1(n_112),
.B2(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_133),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_125),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_143),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_150),
.Y(n_167)
);

AND4x2_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_85),
.C(n_90),
.D(n_100),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_74),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_66),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_73),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_90),
.B1(n_85),
.B2(n_59),
.Y(n_172)
);

NAND4xp75_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_58),
.C(n_59),
.D(n_61),
.Y(n_173)
);

OAI21x1_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_73),
.B(n_71),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_66),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_61),
.C(n_65),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_72),
.B(n_65),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_162),
.C(n_166),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_71),
.A3(n_168),
.B1(n_99),
.B2(n_98),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_109),
.B(n_99),
.C(n_98),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_63),
.B1(n_109),
.B2(n_102),
.C(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_114),
.B(n_118),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_173),
.A3(n_27),
.B1(n_114),
.B2(n_103),
.C1(n_118),
.C2(n_113),
.Y(n_187)
);

AOI211xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_183),
.B(n_182),
.C(n_181),
.Y(n_188)
);

NOR2x1p5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_103),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NAND4xp25_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_103),
.C(n_118),
.D(n_113),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_189),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_191),
.B(n_187),
.C(n_118),
.Y(n_193)
);


endmodule