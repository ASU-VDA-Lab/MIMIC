module fake_jpeg_25880_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_61),
.B1(n_50),
.B2(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_76),
.B1(n_69),
.B2(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_44),
.B1(n_50),
.B2(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_47),
.Y(n_92)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_65),
.B1(n_64),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_55),
.B1(n_60),
.B2(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_75),
.B1(n_86),
.B2(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_93),
.B1(n_101),
.B2(n_68),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_58),
.B1(n_53),
.B2(n_52),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_56),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_100),
.B(n_0),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_0),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_3),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_91),
.B(n_93),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_20),
.B(n_22),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_96),
.B1(n_98),
.B2(n_4),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_4),
.B(n_5),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_26),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_23),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_3),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_104),
.B1(n_6),
.B2(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_104),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_130),
.C(n_134),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_132),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_27),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_29),
.C(n_30),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_131),
.C(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_128),
.B(n_140),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_143),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_137),
.B(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_135),
.C(n_128),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_31),
.C(n_33),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_34),
.CON(n_151),
.SN(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_35),
.Y(n_152)
);


endmodule