module real_jpeg_11631_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g118 ( 
.A(n_0),
.Y(n_118)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_63),
.B1(n_68),
.B2(n_73),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_63),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_274)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_5),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_39),
.B(n_40),
.C(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_50),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_5),
.A2(n_25),
.B1(n_27),
.B2(n_103),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_5),
.A2(n_128),
.B1(n_153),
.B2(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_32),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_105),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_6),
.A2(n_68),
.B1(n_73),
.B2(n_105),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_109),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_109),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_68),
.B1(n_73),
.B2(n_109),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_48),
.B1(n_68),
.B2(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_48),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_12),
.A2(n_25),
.B1(n_27),
.B2(n_52),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_12),
.A2(n_52),
.B1(n_68),
.B2(n_73),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_13),
.A2(n_34),
.B1(n_68),
.B2(n_73),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_13),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_278)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_15),
.A2(n_25),
.B1(n_27),
.B2(n_111),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_68),
.B1(n_73),
.B2(n_111),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_111),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_78),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_19),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_35),
.CI(n_53),
.CON(n_19),
.SN(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_32),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_21),
.A2(n_32),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_21),
.A2(n_32),
.B1(n_136),
.B2(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_21),
.A2(n_33),
.B(n_91),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_21),
.A2(n_32),
.B1(n_88),
.B2(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_22),
.A2(n_89),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_22),
.A2(n_57),
.B(n_274),
.Y(n_273)
);

OA22x2_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_23),
.A2(n_27),
.B(n_171),
.C(n_173),
.Y(n_170)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_25),
.C(n_29),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_25),
.A2(n_27),
.B1(n_71),
.B2(n_74),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_27),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_30),
.B1(n_39),
.B2(n_44),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_29),
.A2(n_44),
.B(n_103),
.Y(n_123)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_30),
.B(n_103),
.CON(n_172),
.SN(n_172)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_33),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_46),
.B(n_49),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_36),
.A2(n_45),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_36),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_36),
.A2(n_49),
.B(n_298),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_47),
.B1(n_50),
.B2(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_37),
.B(n_51),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_37),
.A2(n_50),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_37),
.A2(n_50),
.B1(n_146),
.B2(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_45),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_38)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_62),
.B(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_50),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.C(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_56),
.A2(n_89),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_64),
.A2(n_65),
.B1(n_85),
.B2(n_86),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_82),
.C(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_75),
.B(n_77),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_66),
.B(n_77),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_66),
.A2(n_75),
.B1(n_179),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_66),
.A2(n_75),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_66),
.A2(n_75),
.B1(n_188),
.B2(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_66),
.A2(n_75),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_67),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_67),
.B(n_103),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_SL g74 ( 
.A(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_71),
.B(n_73),
.C(n_103),
.Y(n_195)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_73),
.B(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_77),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_75),
.A2(n_113),
.B(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.C(n_84),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_82),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_82),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_84),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B(n_90),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_302),
.B(n_315),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_283),
.B(n_301),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_258),
.B(n_282),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_162),
.B(n_239),
.C(n_257),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_138),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_99),
.B(n_138),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_115),
.C(n_126),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_100),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_107),
.C(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_103),
.B(n_128),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_110),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_115),
.B(n_126),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_156),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_117),
.A2(n_118),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_118),
.B(n_175),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_134),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_132),
.B1(n_133),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_128),
.A2(n_153),
.B1(n_203),
.B2(n_211),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_128),
.A2(n_153),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_129),
.B(n_221),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_150),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_139),
.B(n_151),
.C(n_161),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_149),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_143),
.B(n_147),
.C(n_149),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_152),
.B(n_157),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_155),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_153),
.A2(n_205),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_159),
.B(n_180),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_234),
.B(n_238),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_189),
.B(n_233),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_184),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_184),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_181),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_176),
.C(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_174),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B(n_180),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_187),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_187),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_228),
.B(n_232),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_217),
.B(n_227),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_206),
.B(n_216),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_201),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_199),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_215),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_223),
.C(n_226),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_256),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_256),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_243),
.C(n_250),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_249),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_246),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_281),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_268),
.B1(n_279),
.B2(n_280),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_280),
.C(n_281),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_264),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_266),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_294),
.B(n_296),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_273),
.C(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_274),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_300),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_300),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_299),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_288),
.C(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_291),
.B(n_292),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_305),
.C(n_309),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_305),
.CI(n_309),
.CON(n_314),
.SN(n_314)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_310),
.Y(n_317)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_314),
.Y(n_319)
);


endmodule