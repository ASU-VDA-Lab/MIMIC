module fake_jpeg_17394_n_218 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_218);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_6),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_45),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_20),
.B1(n_23),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_50),
.B1(n_34),
.B2(n_19),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_35),
.B1(n_20),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_60),
.B1(n_62),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_64),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_38),
.C(n_39),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_75),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_80),
.Y(n_107)
);

NAND2x1_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_38),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_79),
.B1(n_91),
.B2(n_47),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_39),
.B1(n_34),
.B2(n_19),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_89),
.B1(n_92),
.B2(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_26),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_47),
.B1(n_57),
.B2(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_47),
.B1(n_33),
.B2(n_18),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_32),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_2),
.B(n_3),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_33),
.B1(n_18),
.B2(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_89),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_110),
.B1(n_73),
.B2(n_11),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_68),
.B1(n_78),
.B2(n_89),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_114),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_80),
.B(n_16),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_8),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_15),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_125),
.C(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVxp33_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_123),
.B(n_97),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_74),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_68),
.C(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_119),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_85),
.B1(n_78),
.B2(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_82),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_116),
.B(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_10),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_104),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_11),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_102),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_157),
.B(n_153),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_147),
.C(n_142),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_116),
.B(n_103),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_143),
.B(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_111),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_129),
.B1(n_122),
.B2(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_150),
.B(n_156),
.Y(n_185)
);

AOI321xp33_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_172),
.A3(n_168),
.B1(n_167),
.B2(n_164),
.C(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_176),
.C(n_145),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_96),
.B1(n_99),
.B2(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_96),
.B1(n_112),
.B2(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_12),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_12),
.C(n_13),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_159),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_184),
.C(n_188),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_152),
.CI(n_147),
.CON(n_180),
.SN(n_180)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_186),
.B1(n_173),
.B2(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_149),
.C(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_148),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_177),
.C(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_172),
.B1(n_177),
.B2(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_193),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_166),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_181),
.B(n_180),
.C(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_144),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_185),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_179),
.C(n_180),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_191),
.C(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_201),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_200),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_210),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_204),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_198),
.CI(n_199),
.CON(n_213),
.SN(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_214),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_216),
.Y(n_218)
);


endmodule