module fake_jpeg_8809_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx2_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_21),
.B1(n_15),
.B2(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx10_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_14),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_20),
.Y(n_54)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_52),
.B1(n_25),
.B2(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_15),
.B1(n_21),
.B2(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_37),
.B1(n_32),
.B2(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_75),
.B1(n_77),
.B2(n_62),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_38),
.Y(n_65)
);

XNOR2x1_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_13),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_39),
.B1(n_28),
.B2(n_32),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_54),
.B(n_58),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_R g83 ( 
.A(n_65),
.B(n_49),
.Y(n_83)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_65),
.B(n_75),
.C(n_67),
.D(n_66),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_90),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_98),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_63),
.C(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.C(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_77),
.C(n_64),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_86),
.C(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_82),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_49),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_18),
.C(n_16),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_39),
.B1(n_13),
.B2(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_90),
.B1(n_87),
.B2(n_23),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_110),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_95),
.B1(n_80),
.B2(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_91),
.B(n_100),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_0),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_82),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_18),
.B(n_11),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_1),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_1),
.B(n_2),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_103),
.B1(n_108),
.B2(n_111),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.C(n_7),
.Y(n_127)
);

NOR2x1_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_103),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_114),
.B(n_10),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

OAI221xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_120),
.B1(n_6),
.B2(n_5),
.C(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);


endmodule