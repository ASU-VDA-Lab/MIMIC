module fake_jpeg_24996_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_26),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_28),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_35),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_23),
.B1(n_18),
.B2(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_62),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_78),
.Y(n_112)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_65),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_26),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_39),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_28),
.B1(n_31),
.B2(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_25),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_34),
.B1(n_40),
.B2(n_21),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_54),
.B1(n_48),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_64),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_93),
.Y(n_142)
);

OR2x6_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_44),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_56),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_111),
.B1(n_53),
.B2(n_79),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_73),
.C(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_115),
.C(n_37),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_26),
.Y(n_139)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_35),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_34),
.B1(n_40),
.B2(n_36),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_37),
.C(n_49),
.Y(n_115)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_123),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_131),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_63),
.B1(n_40),
.B2(n_34),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_129),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_62),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_32),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_80),
.B1(n_36),
.B2(n_34),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_88),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_87),
.B1(n_36),
.B2(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_83),
.B1(n_78),
.B2(n_76),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_141),
.B(n_99),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_28),
.B(n_16),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_109),
.C(n_115),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_148),
.C(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_95),
.C(n_92),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_158),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_107),
.B(n_93),
.C(n_106),
.D(n_89),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_139),
.C(n_129),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_155),
.B(n_157),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_89),
.B(n_90),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_119),
.C(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_111),
.B1(n_103),
.B2(n_104),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_156),
.B1(n_170),
.B2(n_160),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_108),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_104),
.B1(n_82),
.B2(n_17),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_35),
.B1(n_20),
.B2(n_17),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_110),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_37),
.C(n_75),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_37),
.C(n_53),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_136),
.B1(n_141),
.B2(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_152),
.B1(n_29),
.B2(n_19),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_192),
.C(n_147),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_110),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_184),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_104),
.B(n_124),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_189),
.B(n_35),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_68),
.B1(n_32),
.B2(n_37),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_32),
.B1(n_37),
.B2(n_29),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_37),
.B1(n_29),
.B2(n_35),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_37),
.C(n_35),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_145),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_204),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_184),
.A2(n_174),
.B1(n_183),
.B2(n_176),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_202),
.B1(n_208),
.B2(n_210),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_148),
.B1(n_149),
.B2(n_172),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_163),
.C(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_192),
.C(n_19),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_211),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_20),
.B(n_17),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_214),
.B(n_215),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_20),
.B1(n_19),
.B2(n_3),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_188),
.B1(n_190),
.B2(n_178),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_181),
.B(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_181),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_35),
.C(n_2),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_229),
.B(n_230),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_209),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_1),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_1),
.C(n_2),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_2),
.B(n_3),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_3),
.B(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_199),
.B1(n_211),
.B2(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_221),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_208),
.B1(n_213),
.B2(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_206),
.B1(n_204),
.B2(n_6),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_4),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_224),
.C(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_228),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_216),
.B(n_6),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_238),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_5),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_252),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_5),
.B(n_6),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_242),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_7),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_259),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_233),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_8),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_243),
.C(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_264),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_244),
.B(n_9),
.C(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_R g267 ( 
.A(n_263),
.B(n_8),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_254),
.B(n_256),
.C(n_10),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_267),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_13),
.C2(n_14),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_268),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_260),
.B(n_14),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.C(n_15),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_15),
.Y(n_272)
);


endmodule