module fake_jpeg_15379_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_21),
.Y(n_56)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_60),
.B1(n_72),
.B2(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_55),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_70),
.B1(n_33),
.B2(n_34),
.Y(n_96)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_18),
.B1(n_33),
.B2(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_43),
.B1(n_18),
.B2(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_86),
.B1(n_99),
.B2(n_29),
.Y(n_115)
);

OR2x4_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_18),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_46),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_42),
.B(n_21),
.C(n_24),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_81),
.B(n_92),
.C(n_28),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_41),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_97),
.C(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_96),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_84),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_42),
.B(n_31),
.C(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_27),
.B1(n_31),
.B2(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_34),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_34),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_25),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_26),
.B(n_30),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_41),
.C(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_38),
.B1(n_44),
.B2(n_39),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_62),
.B1(n_55),
.B2(n_47),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_57),
.B1(n_63),
.B2(n_25),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_123),
.B1(n_75),
.B2(n_87),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_115),
.B1(n_122),
.B2(n_99),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_114),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_130),
.B1(n_131),
.B2(n_80),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_126),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_74),
.B1(n_92),
.B2(n_102),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_77),
.B1(n_75),
.B2(n_80),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_127),
.B(n_77),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_124),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_85),
.B1(n_82),
.B2(n_100),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_41),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_38),
.B1(n_36),
.B2(n_39),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_29),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_46),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_121),
.C(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_25),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_17),
.B(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_28),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_28),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_44),
.B1(n_38),
.B2(n_67),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_67),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_138),
.B1(n_142),
.B2(n_156),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_155),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_107),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_148),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_154),
.C(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_151),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_101),
.B1(n_84),
.B2(n_85),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_41),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_41),
.B(n_89),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_44),
.C(n_52),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_112),
.CI(n_110),
.CON(n_160),
.SN(n_160)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_166),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_120),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_165),
.C(n_173),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_119),
.B1(n_127),
.B2(n_107),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_139),
.B1(n_135),
.B2(n_157),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_184),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_114),
.C(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2x1_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_117),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_137),
.B(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_106),
.B1(n_117),
.B2(n_115),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_124),
.B1(n_155),
.B2(n_111),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_105),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_126),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_208),
.B1(n_176),
.B2(n_177),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_133),
.B1(n_152),
.B2(n_136),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_195),
.A2(n_207),
.B1(n_52),
.B2(n_83),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_185),
.B(n_160),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_165),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_104),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_211),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_156),
.B1(n_142),
.B2(n_138),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_179),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_206),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_175),
.B1(n_164),
.B2(n_171),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_146),
.B1(n_134),
.B2(n_159),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_159),
.B1(n_134),
.B2(n_122),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_83),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_113),
.B(n_128),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_215),
.B(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_160),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.C(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_167),
.C(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_202),
.B1(n_213),
.B2(n_199),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_208),
.B1(n_199),
.B2(n_213),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_174),
.C(n_172),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_231),
.C(n_238),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_232),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_177),
.B(n_172),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_230),
.A2(n_233),
.B(n_193),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_130),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_83),
.B(n_111),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_30),
.C(n_17),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_240),
.B(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_30),
.B1(n_17),
.B2(n_2),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_258),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_206),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_209),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_216),
.C(n_227),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_242),
.C(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_192),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_187),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_217),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_230),
.B(n_233),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_266),
.C(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_13),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_235),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_219),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_278),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_276),
.Y(n_292)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_273),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_274),
.C(n_250),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_30),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_8),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_256),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_16),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_291),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_247),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_287),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_242),
.C(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_266),
.C(n_264),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_272),
.B1(n_265),
.B2(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_244),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_267),
.A2(n_241),
.B1(n_255),
.B2(n_253),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_16),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_297),
.B(n_9),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_12),
.B(n_11),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_301),
.C(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_13),
.C(n_12),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_11),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_310),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_0),
.B(n_1),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_311),
.B(n_5),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_2),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_2),
.C(n_3),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_294),
.B1(n_283),
.B2(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_315),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_286),
.B(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_316),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_3),
.C(n_4),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_321),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_5),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_6),
.B(n_323),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_5),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_6),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_318),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_326),
.B(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_6),
.B(n_312),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_322),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_316),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_333),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_336),
.A2(n_337),
.B(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_339),
.B(n_340),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_334),
.CI(n_338),
.CON(n_344),
.SN(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_336),
.Y(n_345)
);


endmodule