module fake_jpeg_7733_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_28),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_40),
.C(n_35),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_47),
.B(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_52),
.B1(n_36),
.B2(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_55),
.B1(n_49),
.B2(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_89),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_61),
.C(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_55),
.B1(n_52),
.B2(n_43),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_52),
.B1(n_43),
.B2(n_17),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_17),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_72),
.B1(n_70),
.B2(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_68),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_100),
.C(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_67),
.B1(n_60),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_102),
.B1(n_108),
.B2(n_82),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_61),
.C(n_69),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_66),
.B(n_73),
.C(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_40),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_35),
.B1(n_41),
.B2(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_117),
.B1(n_125),
.B2(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_87),
.B(n_77),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_77),
.B1(n_87),
.B2(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_104),
.B1(n_94),
.B2(n_101),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_83),
.C(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_81),
.C(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_93),
.C(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_98),
.B1(n_109),
.B2(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_136),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_124),
.B(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_132),
.B1(n_119),
.B2(n_35),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_97),
.B1(n_96),
.B2(n_104),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_94),
.B(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_103),
.B1(n_93),
.B2(n_41),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_1),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_133),
.B1(n_127),
.B2(n_132),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_147),
.B(n_133),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_120),
.C(n_121),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_146),
.C(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_143),
.B1(n_2),
.B2(n_5),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_50),
.B1(n_14),
.B2(n_13),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_14),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_18),
.C(n_12),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_12),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_137),
.B(n_5),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_154),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.C(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_156),
.Y(n_163)
);

XOR2x2_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_18),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_2),
.B(n_6),
.C(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_6),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_149),
.C(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_143),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_142),
.B(n_157),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_167),
.B(n_168),
.Y(n_171)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_157),
.A3(n_8),
.B(n_10),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_157),
.B(n_8),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_170),
.B(n_163),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_7),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_174),
.B(n_11),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_171),
.B(n_10),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);


endmodule