module real_jpeg_10056_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_66),
.B1(n_69),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_74),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_11),
.B(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_3),
.A2(n_36),
.B1(n_66),
.B2(n_69),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_66),
.B1(n_69),
.B2(n_82),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_43),
.B1(n_66),
.B2(n_69),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_101),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_11),
.A2(n_51),
.B(n_84),
.C(n_152),
.D(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_51),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_49),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_70),
.B(n_167),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_11),
.A2(n_31),
.B(n_45),
.C(n_53),
.D(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_31),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_66),
.B1(n_69),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_15),
.A2(n_66),
.B1(n_69),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_16),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_16),
.A2(n_29),
.B1(n_50),
.B2(n_51),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_29),
.B1(n_66),
.B2(n_69),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_76),
.C(n_91),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_22),
.B(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_25),
.A2(n_30),
.B1(n_38),
.B2(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_30),
.B(n_33),
.C(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_33),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_33),
.B(n_60),
.C(n_61),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_30),
.Y(n_101)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_35),
.B(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_37),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_56),
.C(n_57),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_52),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_44),
.B1(n_55),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_46),
.B(n_51),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_48),
.A2(n_50),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_85),
.B(n_87),
.C(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_85),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_55),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_55),
.A2(n_104),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_60),
.B(n_90),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_60),
.B(n_75),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_71),
.B1(n_72),
.B2(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_69),
.B1(n_85),
.B2(n_86),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_87),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_69),
.B(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_69),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_75),
.B1(n_78),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_70),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_71),
.A2(n_72),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_71),
.B(n_168),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_72),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_75),
.A2(n_173),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_75),
.A2(n_181),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_91),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_80),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_83),
.A2(n_90),
.B1(n_164),
.B2(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_83),
.A2(n_195),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_96),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_90),
.A2(n_94),
.B(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_102),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_93),
.B1(n_102),
.B2(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_126),
.B2(n_127),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_145),
.B(n_227),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_143),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_131),
.B(n_143),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_138),
.A2(n_139),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_141),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_221),
.B(n_226),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_208),
.B(n_220),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_189),
.B(n_207),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_169),
.B(n_188),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_177),
.B(n_187),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_175),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B(n_186),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_191),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_200),
.B2(n_206),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_199),
.C(n_206),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_210),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_216),
.C(n_218),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_212),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);


endmodule