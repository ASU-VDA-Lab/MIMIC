module real_jpeg_24676_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_16;

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_17),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_2),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_16),
.B1(n_17),
.B2(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_4),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_4),
.A2(n_19),
.B1(n_31),
.B2(n_32),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_8),
.A2(n_16),
.B1(n_17),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_66),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_48),
.B(n_65),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_27),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_13),
.B(n_27),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_17),
.B1(n_38),
.B2(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_16),
.B(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_53),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_28),
.B(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_40),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_31),
.A2(n_32),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_34),
.B(n_40),
.C(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_55),
.B(n_64),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_87),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_81),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);


endmodule