module fake_aes_942_n_1058 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1058);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1058;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_844;
wire n_769;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_1041;
wire n_578;
wire n_926;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_947;
wire n_924;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_L g272 ( .A(n_261), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_146), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_158), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_92), .Y(n_275) );
CKINVDCx16_ASAP7_75t_R g276 ( .A(n_76), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_207), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_235), .Y(n_278) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_270), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_89), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_262), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_91), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_94), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_201), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_78), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_108), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_40), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_18), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_147), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_30), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_156), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_109), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_47), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_221), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_113), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g299 ( .A(n_155), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_31), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_224), .Y(n_301) );
INVxp33_ASAP7_75t_SL g302 ( .A(n_80), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_119), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_97), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_100), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_254), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_233), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_118), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_87), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_126), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_116), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_10), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_122), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_101), .Y(n_315) );
INVxp33_ASAP7_75t_SL g316 ( .A(n_6), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_148), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_171), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_176), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_197), .Y(n_320) );
INVxp33_ASAP7_75t_SL g321 ( .A(n_195), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_179), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_34), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_178), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_59), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_162), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_43), .Y(n_327) );
CKINVDCx14_ASAP7_75t_R g328 ( .A(n_213), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_41), .Y(n_329) );
CKINVDCx14_ASAP7_75t_R g330 ( .A(n_5), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_182), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_68), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_79), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_130), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_75), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_105), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_127), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_173), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_164), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_65), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_9), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_165), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_227), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_264), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_185), .Y(n_345) );
INVxp33_ASAP7_75t_L g346 ( .A(n_106), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_211), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_198), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_2), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_45), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_47), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_175), .Y(n_352) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_225), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_192), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_238), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_229), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_99), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_177), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_114), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_58), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_237), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_58), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_76), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_42), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_120), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_22), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_160), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_104), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_246), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_216), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_13), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_24), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_186), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_36), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_93), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_250), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_268), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_84), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_96), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_149), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_154), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_95), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_141), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_188), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_204), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_180), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_121), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_222), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_257), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_258), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_60), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_71), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_172), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_25), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_152), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_65), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_200), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_196), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_137), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_144), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_153), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_19), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_45), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_193), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_23), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_271), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_218), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_161), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_90), .Y(n_410) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_157), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_62), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_269), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_187), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_136), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_85), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_239), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_255), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_260), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_212), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_46), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_371), .B(n_0), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_346), .B(n_0), .Y(n_423) );
OA21x2_ASAP7_75t_L g424 ( .A1(n_304), .A2(n_83), .B(n_82), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_330), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_307), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_299), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_307), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_330), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_371), .B(n_1), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_305), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_307), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_307), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_305), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_361), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_385), .B(n_1), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_280), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_385), .B(n_2), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_307), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_280), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_346), .B(n_3), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_285), .B(n_4), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_361), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_291), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_287), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_395), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_291), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
NOR2xp33_ASAP7_75t_R g452 ( .A(n_328), .B(n_86), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_297), .B(n_4), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_360), .B(n_5), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_388), .B(n_6), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_295), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_295), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_287), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_352), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_446), .B(n_353), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_431), .B(n_322), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_429), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_431), .B(n_322), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_425), .A2(n_430), .B1(n_458), .B2(n_446), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_458), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
BUFx10_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_431), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_422), .A2(n_333), .B1(n_403), .B2(n_276), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
NAND2xp33_ASAP7_75t_SL g471 ( .A(n_430), .B(n_309), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_439), .B(n_289), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_439), .B(n_387), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_431), .B(n_290), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_422), .A2(n_340), .B1(n_349), .B2(n_300), .Y(n_476) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_437), .B(n_401), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_437), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_445), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_437), .B(n_328), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_427), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_429), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_437), .B(n_401), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
NOR2xp33_ASAP7_75t_SL g486 ( .A(n_428), .B(n_389), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_426), .B(n_411), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_432), .B(n_398), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_429), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_442), .A2(n_296), .B1(n_313), .B2(n_293), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_442), .A2(n_325), .B1(n_329), .B2(n_323), .Y(n_493) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_445), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_424), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_443), .B(n_332), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_424), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_424), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_466), .B(n_452), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_497), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_472), .A2(n_459), .B1(n_423), .B2(n_453), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_466), .A2(n_435), .B1(n_441), .B2(n_438), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_466), .A2(n_435), .B1(n_441), .B2(n_438), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_484), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_472), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_484), .B(n_452), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_473), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_487), .B(n_443), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_484), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_497), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_488), .B(n_453), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_472), .Y(n_514) );
NOR3xp33_ASAP7_75t_SL g515 ( .A(n_469), .B(n_340), .C(n_300), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_496), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_475), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_489), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_497), .B(n_454), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_480), .B(n_454), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_475), .A2(n_438), .B1(n_456), .B2(n_441), .Y(n_523) );
AND2x6_ASAP7_75t_L g524 ( .A(n_480), .B(n_275), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_472), .B(n_455), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_497), .B(n_455), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_467), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_477), .B(n_417), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_468), .B(n_272), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_477), .B(n_423), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_475), .A2(n_456), .B1(n_441), .B2(n_449), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_475), .A2(n_316), .B1(n_302), .B2(n_309), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_460), .B(n_349), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_496), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_489), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_478), .B(n_277), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_496), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_475), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g540 ( .A1(n_464), .A2(n_316), .B1(n_302), .B2(n_344), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_477), .B(n_321), .Y(n_541) );
AND3x1_ASAP7_75t_SL g542 ( .A(n_476), .B(n_341), .C(n_335), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_474), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_499), .B(n_278), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_461), .B(n_344), .Y(n_545) );
NOR2x2_ASAP7_75t_L g546 ( .A(n_471), .B(n_369), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_461), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_461), .A2(n_441), .B1(n_456), .B2(n_449), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_461), .B(n_283), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_499), .B(n_282), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_479), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_463), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
INVx8_ASAP7_75t_L g555 ( .A(n_463), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_467), .B(n_351), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_463), .B(n_483), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_463), .B(n_369), .Y(n_560) );
NOR2x2_ASAP7_75t_L g561 ( .A(n_467), .B(n_378), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_483), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_483), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_467), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_481), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_483), .B(n_283), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_481), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_539), .A2(n_378), .B1(n_418), .B2(n_492), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_539), .A2(n_418), .B1(n_493), .B2(n_321), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_551), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_506), .B(n_351), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_539), .A2(n_411), .B1(n_498), .B2(n_372), .Y(n_573) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_539), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_521), .B(n_372), .Y(n_576) );
BUFx4f_ASAP7_75t_SL g577 ( .A(n_545), .Y(n_577) );
CKINVDCx8_ASAP7_75t_R g578 ( .A(n_545), .Y(n_578) );
O2A1O1Ixp5_ASAP7_75t_L g579 ( .A1(n_500), .A2(n_274), .B(n_279), .C(n_273), .Y(n_579) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_514), .B(n_498), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_505), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_525), .A2(n_498), .B1(n_312), .B2(n_318), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_544), .A2(n_498), .B(n_491), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_498), .B1(n_312), .B2(n_318), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_509), .B(n_367), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_540), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_527), .B(n_421), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_526), .A2(n_324), .B1(n_337), .B2(n_301), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_513), .B(n_327), .Y(n_592) );
O2A1O1Ixp5_ASAP7_75t_L g593 ( .A1(n_500), .A2(n_342), .B(n_347), .C(n_331), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_534), .B(n_350), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_563), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_560), .B(n_436), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_511), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_533), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_560), .A2(n_451), .B1(n_450), .B2(n_448), .C1(n_447), .C2(n_444), .Y(n_599) );
OAI22xp5_ASAP7_75t_SL g600 ( .A1(n_556), .A2(n_502), .B1(n_510), .B2(n_541), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_515), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_511), .Y(n_602) );
BUFx4f_ASAP7_75t_SL g603 ( .A(n_564), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_547), .Y(n_605) );
NOR2xp67_ASAP7_75t_L g606 ( .A(n_501), .B(n_456), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_SL g607 ( .A1(n_558), .A2(n_457), .B(n_444), .C(n_447), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_557), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_543), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_507), .A2(n_337), .B1(n_345), .B2(n_324), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_516), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_522), .A2(n_363), .B(n_365), .C(n_364), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_541), .B(n_373), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_558), .A2(n_457), .B(n_392), .C(n_393), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_550), .A2(n_490), .B(n_485), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_512), .A2(n_394), .B1(n_396), .B2(n_370), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_529), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_531), .B(n_375), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_552), .A2(n_420), .B1(n_404), .B2(n_412), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_555), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_523), .B(n_397), .Y(n_622) );
OR2x6_ASAP7_75t_SL g623 ( .A(n_561), .B(n_356), .Y(n_623) );
INVx3_ASAP7_75t_SL g624 ( .A(n_546), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_553), .A2(n_448), .B(n_450), .C(n_436), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_523), .B(n_451), .Y(n_626) );
INVx4_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_516), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g629 ( .A1(n_532), .A2(n_357), .B1(n_382), .B2(n_356), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_548), .A2(n_503), .B(n_504), .C(n_532), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_549), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_566), .A2(n_377), .B(n_408), .C(n_359), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_508), .B(n_357), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_524), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_542), .A2(n_286), .B1(n_288), .B2(n_284), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_535), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_524), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_548), .A2(n_362), .B1(n_419), .B2(n_292), .C1(n_294), .C2(n_298), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_530), .A2(n_306), .B(n_303), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_518), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_503), .B(n_384), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_519), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_520), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_524), .Y(n_644) );
AND3x1_ASAP7_75t_SL g645 ( .A(n_542), .B(n_310), .C(n_308), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_530), .A2(n_314), .B1(n_315), .B2(n_311), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_536), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_528), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_537), .A2(n_320), .B(n_326), .C(n_319), .Y(n_649) );
INVx3_ASAP7_75t_L g650 ( .A(n_535), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_565), .A2(n_336), .B(n_339), .C(n_334), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_567), .Y(n_652) );
OR2x6_ASAP7_75t_L g653 ( .A(n_535), .B(n_538), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_538), .Y(n_654) );
BUFx12f_ASAP7_75t_L g655 ( .A(n_538), .Y(n_655) );
INVx5_ASAP7_75t_L g656 ( .A(n_538), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_559), .B(n_343), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_571), .B(n_559), .Y(n_658) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_585), .A2(n_559), .B(n_410), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_653), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_579), .A2(n_354), .B(n_348), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_572), .B(n_7), .Y(n_662) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_650), .A2(n_559), .B(n_410), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_627), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_603), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_655), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_593), .A2(n_366), .B(n_355), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_627), .B(n_281), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_608), .B(n_368), .Y(n_669) );
AO21x2_ASAP7_75t_L g670 ( .A1(n_607), .A2(n_376), .B(n_374), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_592), .B(n_618), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_624), .Y(n_672) );
OAI21x1_ASAP7_75t_L g673 ( .A1(n_650), .A2(n_416), .B(n_358), .Y(n_673) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_621), .B(n_281), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_599), .B(n_379), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_596), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_621), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_626), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_626), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_653), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_581), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_600), .B(n_380), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_613), .B(n_619), .Y(n_683) );
BUFx3_ASAP7_75t_L g684 ( .A(n_574), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_625), .Y(n_685) );
AO32x2_ASAP7_75t_L g686 ( .A1(n_600), .A2(n_440), .A3(n_434), .B1(n_433), .B2(n_427), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_653), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_577), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_614), .A2(n_383), .B(n_381), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_622), .A2(n_390), .B1(n_391), .B2(n_386), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_590), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_652), .A2(n_400), .B(n_399), .Y(n_692) );
OR2x6_ASAP7_75t_L g693 ( .A(n_568), .B(n_402), .Y(n_693) );
OAI21x1_ASAP7_75t_L g694 ( .A1(n_615), .A2(n_407), .B(n_405), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_575), .B(n_409), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_574), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_639), .A2(n_414), .B(n_413), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_594), .A2(n_415), .B1(n_317), .B2(n_338), .C(n_440), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_622), .A2(n_338), .B1(n_317), .B2(n_433), .Y(n_699) );
BUFx4f_ASAP7_75t_L g700 ( .A(n_580), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_609), .Y(n_701) );
INVx6_ASAP7_75t_L g702 ( .A(n_656), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_612), .A2(n_482), .B(n_494), .C(n_462), .Y(n_703) );
OR2x6_ASAP7_75t_L g704 ( .A(n_569), .B(n_7), .Y(n_704) );
OA21x2_ASAP7_75t_L g705 ( .A1(n_649), .A2(n_482), .B(n_462), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_575), .B(n_8), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_586), .Y(n_707) );
AO21x2_ASAP7_75t_L g708 ( .A1(n_635), .A2(n_494), .B(n_482), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_595), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_588), .A2(n_494), .B1(n_9), .B2(n_10), .C(n_11), .Y(n_710) );
OAI21x1_ASAP7_75t_L g711 ( .A1(n_640), .A2(n_98), .B(n_88), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_604), .Y(n_712) );
OAI21x1_ASAP7_75t_L g713 ( .A1(n_642), .A2(n_103), .B(n_102), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_631), .B(n_8), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g715 ( .A(n_656), .B(n_11), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_632), .A2(n_12), .B1(n_13), .B2(n_14), .C(n_15), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_578), .B(n_12), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_617), .Y(n_718) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_601), .B(n_14), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_643), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_656), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_582), .Y(n_722) );
OAI21x1_ASAP7_75t_L g723 ( .A1(n_570), .A2(n_110), .B(n_107), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_635), .B(n_15), .C(n_16), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_647), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_623), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_605), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_634), .B(n_17), .Y(n_728) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_657), .A2(n_112), .B(n_111), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_598), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_730) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_606), .A2(n_117), .B(n_115), .Y(n_731) );
OA21x2_ASAP7_75t_L g732 ( .A1(n_648), .A2(n_124), .B(n_123), .Y(n_732) );
AO21x2_ASAP7_75t_L g733 ( .A1(n_606), .A2(n_128), .B(n_125), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_620), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_583), .A2(n_131), .B(n_129), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_582), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_576), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_629), .Y(n_738) );
OAI21x1_ASAP7_75t_L g739 ( .A1(n_597), .A2(n_133), .B(n_132), .Y(n_739) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_630), .A2(n_135), .B(n_134), .Y(n_740) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_611), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_616), .B(n_20), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_637), .B(n_21), .Y(n_743) );
AO31x2_ASAP7_75t_L g744 ( .A1(n_573), .A2(n_22), .A3(n_23), .B(n_24), .Y(n_744) );
OA21x2_ASAP7_75t_L g745 ( .A1(n_646), .A2(n_139), .B(n_138), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_644), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_651), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_641), .B(n_25), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_602), .A2(n_142), .B(n_140), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_638), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_750) );
AO21x2_ASAP7_75t_L g751 ( .A1(n_584), .A2(n_145), .B(n_143), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_589), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_610), .B(n_29), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_611), .Y(n_754) );
AO21x2_ASAP7_75t_L g755 ( .A1(n_587), .A2(n_151), .B(n_150), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_645), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_616), .B(n_29), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_633), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_591), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_671), .A2(n_654), .B1(n_636), .B2(n_628), .C(n_37), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_701), .Y(n_761) );
OA21x2_ASAP7_75t_L g762 ( .A1(n_659), .A2(n_654), .B(n_636), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_704), .A2(n_693), .B1(n_690), .B2(n_700), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_701), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_683), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_37), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_704), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_734), .A2(n_43), .B1(n_44), .B2(n_46), .C(n_48), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_676), .B(n_44), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_693), .B(n_48), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_693), .B(n_49), .Y(n_770) );
INVx4_ASAP7_75t_L g771 ( .A(n_664), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_690), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_772) );
INVx2_ASAP7_75t_SL g773 ( .A(n_666), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_681), .B(n_52), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_750), .A2(n_53), .B(n_54), .C(n_55), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_738), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_682), .A2(n_56), .B1(n_57), .B2(n_59), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_682), .A2(n_56), .B1(n_61), .B2(n_62), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_718), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_756), .A2(n_63), .B1(n_64), .B2(n_66), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_753), .A2(n_756), .B1(n_759), .B2(n_730), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_681), .Y(n_782) );
AO21x2_ASAP7_75t_L g783 ( .A1(n_703), .A2(n_203), .B(n_266), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_742), .A2(n_67), .B1(n_69), .B2(n_70), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_737), .B(n_70), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_714), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_663), .A2(n_205), .B(n_265), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_718), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_726), .A2(n_72), .B1(n_74), .B2(n_75), .C(n_77), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_664), .B(n_700), .Y(n_790) );
AND2x4_ASAP7_75t_L g791 ( .A(n_678), .B(n_679), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_675), .B(n_74), .Y(n_792) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_747), .A2(n_77), .B(n_78), .C(n_79), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_726), .A2(n_80), .B1(n_81), .B2(n_159), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_662), .B(n_81), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_707), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_709), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_717), .A2(n_163), .B1(n_166), .B2(n_167), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_712), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_669), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_691), .B(n_174), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_727), .B(n_263), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_728), .A2(n_181), .B1(n_183), .B2(n_184), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_727), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_706), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_720), .B(n_194), .Y(n_806) );
BUFx12f_ASAP7_75t_L g807 ( .A(n_665), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_740), .A2(n_202), .B(n_206), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_717), .B(n_208), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_685), .A2(n_209), .B(n_210), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_740), .A2(n_214), .B(n_215), .Y(n_811) );
NOR2xp67_ASAP7_75t_L g812 ( .A(n_688), .B(n_217), .Y(n_812) );
BUFx6f_ASAP7_75t_SL g813 ( .A(n_743), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_757), .A2(n_219), .B1(n_220), .B2(n_223), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_743), .A2(n_226), .B1(n_228), .B2(n_230), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_716), .A2(n_231), .B1(n_232), .B2(n_234), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_677), .B(n_240), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_677), .A2(n_241), .B1(n_243), .B2(n_244), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_658), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_692), .B(n_245), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_715), .A2(n_247), .B1(n_248), .B2(n_249), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_715), .A2(n_251), .B1(n_252), .B2(n_253), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_748), .A2(n_256), .B1(n_695), .B2(n_724), .Y(n_823) );
OR2x6_ASAP7_75t_L g824 ( .A(n_668), .B(n_702), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_744), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_752), .A2(n_710), .B1(n_719), .B2(n_689), .Y(n_826) );
INVx1_ASAP7_75t_SL g827 ( .A(n_702), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_673), .Y(n_828) );
INVx2_ASAP7_75t_SL g829 ( .A(n_702), .Y(n_829) );
OAI211xp5_ASAP7_75t_SL g830 ( .A1(n_758), .A2(n_698), .B(n_699), .C(n_725), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_668), .A2(n_674), .B1(n_725), .B2(n_746), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_L g832 ( .A1(n_661), .A2(n_667), .B(n_697), .C(n_746), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_684), .B(n_696), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_708), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_674), .A2(n_672), .B1(n_721), .B2(n_745), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_708), .A2(n_687), .B1(n_660), .B2(n_680), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_684), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_660), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_670), .A2(n_751), .B1(n_755), .B2(n_745), .Y(n_839) );
AOI222xp33_ASAP7_75t_L g840 ( .A1(n_722), .A2(n_736), .B1(n_754), .B2(n_729), .C1(n_713), .C2(n_711), .Y(n_840) );
INVx3_ASAP7_75t_L g841 ( .A(n_722), .Y(n_841) );
AO31x2_ASAP7_75t_L g842 ( .A1(n_686), .A2(n_705), .A3(n_732), .B(n_751), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_741), .A2(n_705), .B1(n_732), .B2(n_744), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_694), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_686), .B(n_670), .Y(n_845) );
INVx4_ASAP7_75t_L g846 ( .A(n_741), .Y(n_846) );
INVx3_ASAP7_75t_L g847 ( .A(n_741), .Y(n_847) );
AND2x4_ASAP7_75t_L g848 ( .A(n_791), .B(n_731), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_761), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_764), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_779), .B(n_686), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_788), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_834), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_796), .B(n_733), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_825), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_844), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_797), .B(n_732), .Y(n_857) );
INVx2_ASAP7_75t_SL g858 ( .A(n_771), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_769), .B(n_749), .Y(n_859) );
OAI211xp5_ASAP7_75t_L g860 ( .A1(n_789), .A2(n_739), .B(n_735), .C(n_723), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_763), .B(n_799), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_804), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_828), .Y(n_863) );
INVx2_ASAP7_75t_SL g864 ( .A(n_771), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_819), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_774), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_842), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_782), .Y(n_868) );
INVx3_ASAP7_75t_L g869 ( .A(n_846), .Y(n_869) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_846), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_768), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_785), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_792), .B(n_781), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_770), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_838), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_843), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_837), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_842), .Y(n_878) );
BUFx2_ASAP7_75t_L g879 ( .A(n_847), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_766), .B(n_795), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_762), .Y(n_881) );
INVx3_ASAP7_75t_L g882 ( .A(n_790), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_762), .Y(n_883) );
OR2x6_ASAP7_75t_L g884 ( .A(n_790), .B(n_803), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_772), .Y(n_885) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_787), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_806), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_826), .B(n_784), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_812), .Y(n_889) );
OR2x2_ASAP7_75t_L g890 ( .A(n_824), .B(n_827), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_824), .B(n_827), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_813), .B(n_773), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_775), .Y(n_893) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_833), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_841), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_793), .B(n_778), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_845), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_813), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_829), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_783), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_777), .B(n_809), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_765), .Y(n_902) );
BUFx3_ASAP7_75t_L g903 ( .A(n_841), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_831), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_817), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_776), .B(n_803), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_836), .B(n_802), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_821), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_786), .B(n_794), .Y(n_909) );
BUFx3_ASAP7_75t_L g910 ( .A(n_807), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_821), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_767), .B(n_801), .Y(n_912) );
INVx2_ASAP7_75t_SL g913 ( .A(n_822), .Y(n_913) );
INVxp67_ASAP7_75t_SL g914 ( .A(n_822), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_835), .A2(n_811), .B(n_808), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_780), .B(n_832), .Y(n_916) );
INVx3_ASAP7_75t_L g917 ( .A(n_820), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_760), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_810), .B(n_816), .Y(n_919) );
OAI211xp5_ASAP7_75t_L g920 ( .A1(n_798), .A2(n_830), .B(n_839), .C(n_823), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_818), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_815), .B(n_805), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_868), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_861), .B(n_800), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_873), .B(n_814), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_856), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_897), .B(n_840), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_856), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_888), .A2(n_880), .B1(n_912), .B2(n_901), .Y(n_929) );
AND2x4_ASAP7_75t_L g930 ( .A(n_855), .B(n_848), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_866), .B(n_874), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_865), .B(n_855), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_865), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_877), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_858), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_853), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_862), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_849), .B(n_850), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_875), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_852), .B(n_854), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_906), .A2(n_918), .B1(n_902), .B2(n_909), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_870), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_864), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_882), .Y(n_944) );
AOI33xp33_ASAP7_75t_L g945 ( .A1(n_872), .A2(n_871), .A3(n_898), .B1(n_893), .B2(n_899), .B3(n_889), .Y(n_945) );
INVx4_ASAP7_75t_L g946 ( .A(n_884), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_918), .A2(n_885), .B1(n_916), .B2(n_896), .C(n_906), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_881), .Y(n_948) );
BUFx2_ASAP7_75t_L g949 ( .A(n_884), .Y(n_949) );
BUFx2_ASAP7_75t_L g950 ( .A(n_870), .Y(n_950) );
OR2x2_ASAP7_75t_L g951 ( .A(n_890), .B(n_891), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_851), .B(n_859), .Y(n_952) );
INVx5_ASAP7_75t_L g953 ( .A(n_882), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_883), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_887), .B(n_882), .Y(n_955) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_903), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_848), .B(n_859), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_913), .A2(n_911), .B1(n_908), .B2(n_904), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_908), .A2(n_911), .B1(n_914), .B2(n_919), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_883), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_915), .A2(n_860), .B(n_920), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_863), .Y(n_962) );
INVx3_ASAP7_75t_SL g963 ( .A(n_910), .Y(n_963) );
BUFx2_ASAP7_75t_L g964 ( .A(n_869), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_921), .A2(n_905), .B1(n_922), .B2(n_892), .C(n_907), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_863), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_869), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_952), .B(n_876), .Y(n_968) );
NAND2xp5_ASAP7_75t_SL g969 ( .A(n_945), .B(n_894), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_963), .Y(n_970) );
INVx1_ASAP7_75t_SL g971 ( .A(n_963), .Y(n_971) );
AND2x4_ASAP7_75t_L g972 ( .A(n_930), .B(n_848), .Y(n_972) );
AND2x4_ASAP7_75t_SL g973 ( .A(n_946), .B(n_894), .Y(n_973) );
INVx2_ASAP7_75t_SL g974 ( .A(n_967), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_937), .Y(n_975) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_935), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_939), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_940), .B(n_867), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_948), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_932), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_941), .B(n_879), .Y(n_981) );
NOR2xp67_ASAP7_75t_SL g982 ( .A(n_946), .B(n_894), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_957), .B(n_878), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_923), .Y(n_984) );
BUFx3_ASAP7_75t_L g985 ( .A(n_943), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_957), .B(n_857), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_931), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_941), .B(n_895), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_947), .B(n_895), .Y(n_989) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_945), .B(n_917), .C(n_900), .Y(n_990) );
BUFx2_ASAP7_75t_L g991 ( .A(n_946), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_933), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_929), .B(n_917), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_954), .Y(n_994) );
CKINVDCx11_ASAP7_75t_R g995 ( .A(n_934), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_954), .Y(n_996) );
NAND2x1p5_ASAP7_75t_L g997 ( .A(n_953), .B(n_917), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_964), .Y(n_998) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_956), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_950), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_927), .B(n_886), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_930), .B(n_886), .Y(n_1002) );
INVxp67_ASAP7_75t_L g1003 ( .A(n_992), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_987), .B(n_959), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_986), .B(n_951), .Y(n_1005) );
NOR3xp33_ASAP7_75t_SL g1006 ( .A(n_970), .B(n_965), .C(n_961), .Y(n_1006) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_972), .B(n_949), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_975), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_968), .B(n_959), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_977), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_984), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_980), .B(n_958), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1013 ( .A(n_985), .Y(n_1013) );
AND2x4_ASAP7_75t_SL g1014 ( .A(n_999), .B(n_942), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_976), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1016 ( .A(n_1000), .Y(n_1016) );
AND2x4_ASAP7_75t_SL g1017 ( .A(n_972), .B(n_942), .Y(n_1017) );
INVx1_ASAP7_75t_SL g1018 ( .A(n_970), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_974), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_989), .B(n_925), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_983), .B(n_938), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_998), .B(n_936), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1008), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1010), .Y(n_1024) );
AOI321xp33_ASAP7_75t_L g1025 ( .A1(n_1020), .A2(n_993), .A3(n_988), .B1(n_981), .B2(n_969), .C(n_1001), .Y(n_1025) );
NAND3xp33_ASAP7_75t_L g1026 ( .A(n_1006), .B(n_990), .C(n_995), .Y(n_1026) );
NOR2xp33_ASAP7_75t_L g1027 ( .A(n_1020), .B(n_971), .Y(n_1027) );
NAND2x1_ASAP7_75t_L g1028 ( .A(n_1013), .B(n_982), .Y(n_1028) );
INVx1_ASAP7_75t_SL g1029 ( .A(n_1018), .Y(n_1029) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_1016), .Y(n_1030) );
NAND2xp5_ASAP7_75t_SL g1031 ( .A(n_1013), .B(n_991), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_1004), .A2(n_955), .B1(n_997), .B2(n_924), .C(n_982), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1022), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_1003), .A2(n_997), .B1(n_953), .B2(n_944), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1009), .B(n_978), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_1027), .B(n_1003), .Y(n_1036) );
O2A1O1Ixp5_ASAP7_75t_L g1037 ( .A1(n_1031), .A2(n_1015), .B(n_1016), .C(n_1011), .Y(n_1037) );
INVx1_ASAP7_75t_SL g1038 ( .A(n_1029), .Y(n_1038) );
NAND2xp5_ASAP7_75t_SL g1039 ( .A(n_1031), .B(n_1019), .Y(n_1039) );
INVxp33_ASAP7_75t_L g1040 ( .A(n_1028), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1023), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1035), .B(n_1005), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1040), .B(n_1033), .Y(n_1043) );
AO22x2_ASAP7_75t_L g1044 ( .A1(n_1038), .A2(n_1026), .B1(n_1030), .B2(n_1024), .Y(n_1044) );
OAI21xp5_ASAP7_75t_L g1045 ( .A1(n_1037), .A2(n_1039), .B(n_1040), .Y(n_1045) );
OAI31xp33_ASAP7_75t_SL g1046 ( .A1(n_1039), .A2(n_1034), .A3(n_1032), .B(n_1007), .Y(n_1046) );
AND2x2_ASAP7_75t_SL g1047 ( .A(n_1036), .B(n_1014), .Y(n_1047) );
O2A1O1Ixp5_ASAP7_75t_SL g1048 ( .A1(n_1045), .A2(n_1041), .B(n_1042), .C(n_1012), .Y(n_1048) );
A2O1A1Ixp33_ASAP7_75t_L g1049 ( .A1(n_1046), .A2(n_1025), .B(n_1014), .C(n_1017), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1047), .A2(n_1007), .B1(n_1021), .B2(n_973), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_1050), .A2(n_1044), .B1(n_1047), .B2(n_1043), .Y(n_1051) );
NAND3xp33_ASAP7_75t_SL g1052 ( .A(n_1051), .B(n_1048), .C(n_1049), .Y(n_1052) );
XNOR2xp5_ASAP7_75t_L g1053 ( .A(n_1052), .B(n_1002), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1053), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1054), .Y(n_1055) );
OA21x2_ASAP7_75t_L g1056 ( .A1(n_1055), .A2(n_928), .B(n_926), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_1056), .A2(n_979), .B1(n_996), .B2(n_994), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_1057), .A2(n_960), .B1(n_962), .B2(n_966), .Y(n_1058) );
endmodule