module fake_jpeg_10954_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_50),
.Y(n_89)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_59),
.Y(n_81)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_3),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_60),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_65),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_69),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_24),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_26),
.B1(n_16),
.B2(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_95),
.B1(n_113),
.B2(n_60),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_82),
.B(n_117),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_16),
.B1(n_38),
.B2(n_27),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_74),
.B1(n_58),
.B2(n_12),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_84),
.A2(n_11),
.B1(n_102),
.B2(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_103),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_36),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_108),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_43),
.B(n_20),
.C(n_70),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_110),
.B(n_104),
.C(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_114),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_9),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_52),
.B(n_9),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_57),
.B1(n_65),
.B2(n_67),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_130),
.B1(n_136),
.B2(n_138),
.Y(n_169)
);

NAND2x1_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_71),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_149),
.C(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_142),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_58),
.B1(n_10),
.B2(n_11),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_83),
.A2(n_11),
.B1(n_86),
.B2(n_91),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_115),
.B1(n_97),
.B2(n_99),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_144),
.B1(n_141),
.B2(n_147),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_106),
.B1(n_117),
.B2(n_110),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_148),
.Y(n_177)
);

AOI211xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_87),
.B(n_101),
.C(n_109),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_92),
.C(n_85),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_101),
.B1(n_115),
.B2(n_99),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_146),
.B1(n_127),
.B2(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_89),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_89),
.B(n_97),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_87),
.B(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_157),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_79),
.A2(n_112),
.B(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_93),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_79),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_101),
.B1(n_87),
.B2(n_116),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_178),
.B1(n_129),
.B2(n_154),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_165),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_170),
.B(n_129),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_93),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_109),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_87),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_148),
.C(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_138),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_129),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_130),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_191),
.C(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_193),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_161),
.B1(n_135),
.B2(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_166),
.B(n_177),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_195),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_197),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_152),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_133),
.C(n_145),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_135),
.B1(n_137),
.B2(n_123),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_134),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_139),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_165),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_181),
.B(n_172),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_217),
.B(n_188),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_166),
.B1(n_170),
.B2(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_182),
.B1(n_183),
.B2(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_169),
.B1(n_180),
.B2(n_167),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_198),
.B1(n_203),
.B2(n_194),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_169),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_166),
.C(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_182),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_177),
.C(n_171),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_173),
.B(n_160),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_199),
.Y(n_225)
);

OA21x2_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_206),
.B(n_214),
.Y(n_233)
);

AOI31xp67_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_189),
.A3(n_205),
.B(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

OA21x2_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_217),
.B(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_211),
.B1(n_207),
.B2(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_240),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_239),
.B(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_245),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_246),
.B1(n_237),
.B2(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_208),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_227),
.C(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_215),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_235),
.B(n_237),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_229),
.B(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_244),
.C(n_240),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_236),
.B1(n_238),
.B2(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_254),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_250),
.B(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_228),
.Y(n_261)
);


endmodule