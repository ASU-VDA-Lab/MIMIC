module fake_jpeg_25515_n_98 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_29),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_1),
.Y(n_42)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_20),
.B1(n_19),
.B2(n_13),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_36),
.B1(n_42),
.B2(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_11),
.B1(n_22),
.B2(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_30),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_34),
.C(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_31),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_46),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_28),
.B1(n_27),
.B2(n_34),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_62),
.B1(n_48),
.B2(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_27),
.B1(n_24),
.B2(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_24),
.C(n_7),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_66),
.C(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_46),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_1),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_66),
.C(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_75),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_46),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_45),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_82),
.B1(n_2),
.B2(n_4),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_2),
.C(n_78),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_70),
.B(n_3),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_87),
.C(n_81),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_85),
.C(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_86),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_92),
.Y(n_98)
);


endmodule