module fake_netlist_5_2439_n_116 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_53, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_51, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_3, n_49, n_52, n_6, n_39, n_116);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_51;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_3;
input n_49;
input n_52;
input n_6;
input n_39;

output n_116;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_111;
wire n_108;
wire n_66;
wire n_98;
wire n_60;
wire n_107;
wire n_58;
wire n_69;
wire n_94;
wire n_113;
wire n_105;
wire n_80;
wire n_73;
wire n_92;
wire n_84;
wire n_79;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_59;
wire n_99;
wire n_67;
wire n_76;
wire n_87;
wire n_77;
wire n_102;
wire n_106;
wire n_64;
wire n_81;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_104;
wire n_103;
wire n_56;
wire n_63;
wire n_97;
wire n_88;
wire n_110;

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_23),
.A2(n_44),
.B1(n_54),
.B2(n_4),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_19),
.B(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_13),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_10),
.B1(n_42),
.B2(n_0),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_24),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_37),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_27),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_11),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AND3x2_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_2),
.C(n_6),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_2),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_7),
.B1(n_12),
.B2(n_14),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_16),
.B1(n_20),
.B2(n_29),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_71),
.B(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_63),
.B1(n_76),
.B2(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_68),
.B(n_63),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_61),
.B(n_77),
.Y(n_95)
);

AO31x2_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_56),
.A3(n_59),
.B(n_60),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_73),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_95),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_80),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_90),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_97),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_102),
.Y(n_108)
);

NAND2x1_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_60),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_104),
.B(n_105),
.C(n_103),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_104),
.B(n_74),
.C(n_81),
.Y(n_111)
);

OR5x1_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_64),
.C(n_89),
.D(n_79),
.E(n_74),
.Y(n_112)
);

OAI211xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_79),
.B(n_67),
.C(n_34),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_30),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_113),
.B1(n_36),
.B2(n_39),
.Y(n_115)
);

OA331x2_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_32),
.A3(n_40),
.B1(n_46),
.B2(n_49),
.B3(n_50),
.C1(n_55),
.Y(n_116)
);


endmodule