module fake_netlist_6_3492_n_1611 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1611);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1611;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_43),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_40),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_40),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_42),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_3),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_92),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_1),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_19),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_94),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_45),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_73),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_65),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_78),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_85),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_80),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_21),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_15),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_44),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_57),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_104),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_20),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_71),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_27),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_30),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_11),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_19),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_90),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_98),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_70),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_44),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_55),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_89),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_53),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_83),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_130),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_38),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_95),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_59),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_72),
.Y(n_230)
);

BUFx2_ASAP7_75t_SL g231 ( 
.A(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_22),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_61),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_29),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_34),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_49),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_67),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_7),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_57),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_25),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_84),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_22),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_50),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_3),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_58),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_62),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_102),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_4),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_8),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_36),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_133),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_14),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_53),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_35),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_24),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_49),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_52),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_26),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_142),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_152),
.B(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_143),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_206),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_152),
.B(n_5),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_193),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_149),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_157),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_161),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_162),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_164),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_165),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_147),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_171),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_273),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_202),
.B(n_12),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_273),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_148),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_173),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_155),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_170),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_175),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_192),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_206),
.B(n_12),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_211),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_192),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_176),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_178),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_177),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_222),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_183),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_179),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_208),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_177),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_169),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_177),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_144),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_144),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_154),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_154),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_181),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_158),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_189),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_191),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_247),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_284),
.B(n_247),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_287),
.B(n_203),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_156),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_289),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_289),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_290),
.B(n_203),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_297),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_290),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_293),
.B(n_209),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_209),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_150),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_295),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_150),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_300),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_346),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_300),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_301),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_297),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_151),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_L g414 ( 
.A(n_333),
.B(n_202),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_322),
.B(n_276),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_340),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_347),
.B(n_151),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_286),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_349),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_285),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_365),
.B(n_294),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

BUFx4f_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

BUFx6f_ASAP7_75t_SL g434 ( 
.A(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_303),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_306),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_307),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_361),
.B(n_310),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_350),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx4_ASAP7_75t_SL g451 ( 
.A(n_378),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_377),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

BUFx4f_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_361),
.B(n_314),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_315),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_R g466 ( 
.A(n_401),
.B(n_317),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_405),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_374),
.B(n_320),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_374),
.B(n_311),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_388),
.A2(n_358),
.B1(n_299),
.B2(n_355),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_397),
.B(n_153),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_327),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_388),
.B(n_331),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_406),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_406),
.B(n_336),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_405),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_414),
.A2(n_296),
.B1(n_276),
.B2(n_185),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

BUFx4f_ASAP7_75t_L g488 ( 
.A(n_378),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_378),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_378),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_415),
.B(n_337),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_378),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_369),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_412),
.B(n_185),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_426),
.B(n_342),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_420),
.A2(n_357),
.B1(n_298),
.B2(n_291),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_420),
.A2(n_326),
.B1(n_237),
.B2(n_215),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_369),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_378),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_369),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_369),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_183),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_419),
.B(n_421),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_419),
.B(n_350),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_370),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_L g511 ( 
.A(n_414),
.B(n_197),
.C(n_182),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_389),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_384),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_344),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_389),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_412),
.A2(n_194),
.B1(n_275),
.B2(n_278),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_389),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_359),
.B(n_305),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_397),
.B(n_168),
.C(n_153),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_391),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_359),
.B(n_201),
.C(n_198),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_384),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_391),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_397),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_397),
.A2(n_275),
.B1(n_194),
.B2(n_249),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_360),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_363),
.B(n_325),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_370),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_393),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_363),
.B(n_248),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_396),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_400),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_393),
.B(n_168),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_393),
.A2(n_283),
.B1(n_187),
.B2(n_146),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_363),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_400),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_400),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_400),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_364),
.B(n_204),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_421),
.B(n_345),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_364),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_362),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_364),
.B(n_351),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_393),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_370),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_421),
.B(n_345),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_393),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_393),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_427),
.B(n_328),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_370),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_393),
.B(n_195),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_362),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_362),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_395),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_427),
.B(n_329),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_366),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_370),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_386),
.B(n_183),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_366),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_386),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_508),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_568),
.B(n_395),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_481),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_566),
.B(n_395),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_541),
.B(n_218),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_220),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_479),
.B(n_158),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_489),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_484),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_395),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_481),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_484),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_566),
.B(n_395),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_441),
.B(n_395),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_483),
.A2(n_390),
.B(n_368),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_527),
.B(n_395),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_444),
.A2(n_166),
.B1(n_172),
.B2(n_184),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_466),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_515),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_442),
.B(n_402),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_550),
.A2(n_238),
.B(n_186),
.C(n_205),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_535),
.B(n_196),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_459),
.B(n_402),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_547),
.A2(n_334),
.B1(n_230),
.B2(n_259),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_477),
.B(n_402),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_546),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_550),
.B(n_402),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_551),
.B(n_402),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_551),
.B(n_402),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_556),
.B(n_402),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_428),
.B(n_402),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_444),
.B(n_402),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_473),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_556),
.B(n_402),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_546),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_519),
.B(n_404),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_429),
.B(n_404),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_487),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_435),
.B(n_404),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_531),
.B(n_404),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_478),
.B(n_228),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_404),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_487),
.B(n_351),
.Y(n_619)
);

O2A1O1Ixp5_ASAP7_75t_L g620 ( 
.A1(n_475),
.A2(n_390),
.B(n_366),
.C(n_367),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_475),
.B(n_174),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_485),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_475),
.A2(n_238),
.B1(n_205),
.B2(n_216),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_475),
.B(n_404),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_540),
.A2(n_225),
.B1(n_219),
.B2(n_216),
.C(n_232),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_553),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_507),
.B(n_404),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_522),
.B(n_427),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_437),
.B(n_404),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_437),
.B(n_445),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_553),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_474),
.B(n_390),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_497),
.B(n_219),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_506),
.A2(n_266),
.B(n_246),
.C(n_249),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_473),
.B(n_229),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_548),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_434),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_560),
.A2(n_561),
.B(n_559),
.C(n_500),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_536),
.A2(n_545),
.B1(n_563),
.B2(n_557),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_445),
.B(n_404),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_539),
.A2(n_272),
.B1(n_260),
.B2(n_246),
.Y(n_645)
);

INVxp33_ASAP7_75t_SL g646 ( 
.A(n_540),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_430),
.B(n_234),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_501),
.A2(n_239),
.B1(n_232),
.B2(n_225),
.C(n_255),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_446),
.B(n_404),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_482),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_497),
.B(n_236),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_443),
.B(n_240),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_487),
.B(n_352),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_446),
.B(n_183),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_458),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_447),
.B(n_423),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_447),
.B(n_183),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_539),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_448),
.B(n_423),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_448),
.B(n_423),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_539),
.A2(n_239),
.B1(n_255),
.B2(n_260),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_450),
.B(n_423),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_470),
.B(n_263),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_517),
.A2(n_263),
.B(n_266),
.C(n_272),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_528),
.A2(n_278),
.B(n_262),
.C(n_235),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_450),
.B(n_183),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_485),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_452),
.B(n_188),
.Y(n_669)
);

NAND2x1_ASAP7_75t_L g670 ( 
.A(n_530),
.B(n_360),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_480),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_493),
.B(n_243),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_511),
.B(n_244),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_452),
.B(n_423),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_455),
.B(n_423),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_498),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_455),
.B(n_367),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_456),
.B(n_367),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_456),
.B(n_372),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_434),
.A2(n_224),
.B1(n_199),
.B2(n_207),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_461),
.B(n_372),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_486),
.B(n_188),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_461),
.B(n_188),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_485),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_485),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_465),
.B(n_372),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_564),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_210),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_465),
.B(n_245),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_525),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_509),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_520),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_467),
.B(n_373),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_467),
.B(n_373),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_525),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_468),
.B(n_373),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_468),
.B(n_250),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_509),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_509),
.Y(n_701)
);

INVx8_ASAP7_75t_L g702 ( 
.A(n_434),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_469),
.A2(n_381),
.B(n_375),
.C(n_380),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_434),
.A2(n_200),
.B1(n_190),
.B2(n_262),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_469),
.B(n_375),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_476),
.B(n_268),
.C(n_252),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_525),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_476),
.A2(n_221),
.B1(n_200),
.B2(n_214),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_490),
.B(n_375),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_496),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_496),
.B(n_380),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_549),
.B(n_188),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_509),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_510),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_510),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_509),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_549),
.B(n_188),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_513),
.B(n_516),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_554),
.B(n_180),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_554),
.B(n_212),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_554),
.B(n_270),
.C(n_271),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_513),
.B(n_352),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_586),
.A2(n_457),
.B(n_432),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_582),
.A2(n_457),
.B(n_432),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_592),
.A2(n_457),
.B(n_432),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_596),
.A2(n_457),
.B(n_432),
.Y(n_727)
);

BUFx4f_ASAP7_75t_L g728 ( 
.A(n_635),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_634),
.B(n_509),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_585),
.A2(n_488),
.B(n_516),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_600),
.A2(n_488),
.B(n_518),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_643),
.B(n_558),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_641),
.A2(n_235),
.B(n_233),
.C(n_214),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_710),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_574),
.A2(n_488),
.B(n_518),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_606),
.B(n_521),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_637),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_569),
.B(n_524),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_570),
.B(n_591),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_578),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_619),
.B(n_353),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_595),
.B(n_524),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_601),
.B(n_562),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_658),
.A2(n_530),
.B1(n_562),
.B2(n_529),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_578),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_639),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_617),
.A2(n_530),
.B1(n_562),
.B2(n_529),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_716),
.A2(n_488),
.B(n_471),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_716),
.A2(n_471),
.B(n_436),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_716),
.A2(n_471),
.B(n_436),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_610),
.B(n_565),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_670),
.A2(n_471),
.B(n_436),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_667),
.A2(n_491),
.B(n_436),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_621),
.B(n_353),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_627),
.B(n_438),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_602),
.A2(n_492),
.B(n_491),
.Y(n_756)
);

NOR2x2_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_253),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_633),
.B(n_565),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_578),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_653),
.B(n_558),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_579),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_640),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_611),
.A2(n_538),
.B(n_532),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_598),
.B(n_558),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_612),
.A2(n_492),
.B(n_491),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_647),
.B(n_213),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_615),
.A2(n_494),
.B(n_492),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_590),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_572),
.A2(n_543),
.B1(n_494),
.B2(n_492),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_608),
.B(n_494),
.Y(n_770)
);

BUFx8_ASAP7_75t_L g771 ( 
.A(n_613),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_574),
.A2(n_449),
.B(n_431),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_640),
.B(n_226),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_655),
.B(n_217),
.Y(n_774)
);

AOI21x1_ASAP7_75t_L g775 ( 
.A1(n_611),
.A2(n_433),
.B(n_472),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_588),
.A2(n_587),
.B(n_618),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_704),
.A2(n_227),
.B1(n_552),
.B2(n_533),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_671),
.B(n_223),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_620),
.A2(n_453),
.B(n_431),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_642),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_704),
.A2(n_227),
.B1(n_552),
.B2(n_533),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_652),
.B(n_241),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_575),
.B(n_438),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_631),
.B(n_494),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_575),
.B(n_576),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_668),
.Y(n_786)
);

AO21x1_ASAP7_75t_L g787 ( 
.A1(n_616),
.A2(n_673),
.B(n_622),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_663),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_576),
.B(n_565),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_571),
.B(n_438),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_689),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_616),
.A2(n_463),
.B(n_544),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_SL g793 ( 
.A1(n_625),
.A2(n_534),
.B(n_537),
.C(n_542),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_588),
.A2(n_503),
.B(n_460),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_628),
.A2(n_503),
.B(n_460),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_503),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_638),
.B(n_354),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_593),
.A2(n_537),
.B(n_544),
.C(n_542),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_635),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_607),
.A2(n_632),
.B(n_625),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_603),
.A2(n_433),
.B(n_472),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_665),
.A2(n_664),
.B(n_708),
.C(n_580),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_614),
.A2(n_503),
.B(n_460),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_665),
.A2(n_537),
.B(n_463),
.C(n_439),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_614),
.A2(n_460),
.B(n_495),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_581),
.A2(n_552),
.B1(n_533),
.B2(n_438),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_614),
.A2(n_460),
.B(n_495),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_691),
.B(n_552),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_652),
.B(n_440),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_614),
.A2(n_460),
.B(n_495),
.Y(n_810)
);

BUFx5_ASAP7_75t_L g811 ( 
.A(n_584),
.Y(n_811)
);

BUFx4f_ASAP7_75t_L g812 ( 
.A(n_663),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_699),
.B(n_533),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_599),
.B(n_673),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_623),
.A2(n_495),
.B(n_360),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_699),
.B(n_440),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_SL g817 ( 
.A1(n_649),
.A2(n_526),
.B(n_523),
.C(n_514),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_623),
.A2(n_495),
.B(n_360),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_714),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_631),
.B(n_242),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_629),
.A2(n_454),
.B1(n_505),
.B2(n_504),
.Y(n_821)
);

AO21x1_ASAP7_75t_L g822 ( 
.A1(n_622),
.A2(n_526),
.B(n_523),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_623),
.A2(n_495),
.B(n_360),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_664),
.A2(n_514),
.B(n_512),
.C(n_439),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_684),
.A2(n_454),
.B1(n_505),
.B2(n_504),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_623),
.A2(n_360),
.B(n_505),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_715),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_684),
.A2(n_512),
.B(n_449),
.C(n_453),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_706),
.B(n_258),
.Y(n_829)
);

AO21x1_ASAP7_75t_L g830 ( 
.A1(n_718),
.A2(n_392),
.B(n_399),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_722),
.B(n_505),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_656),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_675),
.A2(n_360),
.B(n_502),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_694),
.B(n_354),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_718),
.B(n_440),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_624),
.B(n_440),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_626),
.A2(n_504),
.B(n_502),
.C(n_464),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_SL g838 ( 
.A1(n_649),
.A2(n_604),
.B(n_603),
.C(n_609),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_577),
.B(n_356),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_648),
.A2(n_504),
.B(n_502),
.C(n_464),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_630),
.A2(n_502),
.B(n_464),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_659),
.Y(n_842)
);

INVx11_ASAP7_75t_L g843 ( 
.A(n_651),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_624),
.B(n_464),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_675),
.A2(n_454),
.B(n_370),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_605),
.A2(n_370),
.B(n_368),
.Y(n_846)
);

NOR2x1_ASAP7_75t_R g847 ( 
.A(n_654),
.B(n_254),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_605),
.A2(n_370),
.B(n_368),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_686),
.B(n_451),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_609),
.A2(n_370),
.B(n_368),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_675),
.B(n_381),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_577),
.B(n_356),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_660),
.A2(n_381),
.B(n_382),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_687),
.B(n_451),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_640),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_719),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_644),
.A2(n_370),
.B(n_371),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_662),
.A2(n_371),
.B(n_376),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_703),
.A2(n_392),
.B(n_409),
.C(n_407),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_672),
.B(n_256),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_674),
.A2(n_371),
.B(n_376),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_676),
.A2(n_371),
.B(n_376),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_679),
.A2(n_385),
.B(n_382),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_SL g864 ( 
.A(n_702),
.B(n_267),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_687),
.B(n_451),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_682),
.A2(n_279),
.B(n_424),
.C(n_410),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_680),
.A2(n_387),
.B(n_392),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_681),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_683),
.A2(n_376),
.B(n_371),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_693),
.B(n_713),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_688),
.A2(n_376),
.B(n_371),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_695),
.A2(n_376),
.B(n_409),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_693),
.B(n_451),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_696),
.A2(n_387),
.B(n_382),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_589),
.B(n_348),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_698),
.A2(n_424),
.B(n_410),
.C(n_413),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_702),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_713),
.B(n_385),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_705),
.A2(n_711),
.B(n_709),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_573),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_675),
.A2(n_700),
.B(n_701),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_654),
.A2(n_407),
.B(n_387),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_583),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_657),
.A2(n_409),
.B(n_398),
.C(n_399),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_700),
.A2(n_385),
.B(n_398),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_700),
.A2(n_398),
.B(n_399),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_650),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_700),
.A2(n_403),
.B(n_424),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_768),
.B(n_855),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_785),
.A2(n_589),
.B1(n_645),
.B2(n_661),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_761),
.B(n_594),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_860),
.A2(n_690),
.B(n_721),
.C(n_661),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_737),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_740),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_748),
.A2(n_701),
.B(n_702),
.Y(n_895)
);

NOR2x1_ASAP7_75t_SL g896 ( 
.A(n_740),
.B(n_701),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_868),
.B(n_645),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_797),
.B(n_741),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_832),
.B(n_677),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_782),
.A2(n_666),
.B(n_685),
.C(n_669),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_746),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_749),
.A2(n_701),
.B(n_720),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_875),
.A2(n_719),
.B1(n_697),
.B2(n_678),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_766),
.A2(n_707),
.B1(n_692),
.B2(n_723),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_740),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_796),
.A2(n_636),
.B(n_669),
.C(n_685),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_780),
.Y(n_907)
);

CKINVDCx8_ASAP7_75t_R g908 ( 
.A(n_855),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_786),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_776),
.A2(n_717),
.B(n_712),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_819),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_791),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_812),
.B(n_281),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_827),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_739),
.A2(n_280),
.B1(n_265),
.B2(n_269),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_809),
.A2(n_261),
.B(n_274),
.C(n_277),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_855),
.Y(n_917)
);

AOI221xp5_ASAP7_75t_L g918 ( 
.A1(n_834),
.A2(n_417),
.B1(n_413),
.B2(n_410),
.C(n_422),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_771),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_842),
.B(n_417),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_754),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_SL g922 ( 
.A1(n_770),
.A2(n_410),
.B(n_417),
.C(n_413),
.Y(n_922)
);

INVx3_ASAP7_75t_SL g923 ( 
.A(n_757),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_750),
.A2(n_417),
.B(n_413),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_788),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_738),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_864),
.B(n_64),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_742),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_880),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_745),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_725),
.A2(n_879),
.B(n_736),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_745),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_732),
.A2(n_410),
.B(n_413),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_879),
.A2(n_422),
.B(n_418),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_852),
.B(n_422),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_774),
.B(n_13),
.C(n_14),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_831),
.A2(n_422),
.B(n_418),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_883),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_759),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_733),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_783),
.B(n_422),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_759),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_789),
.B(n_422),
.C(n_418),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_808),
.A2(n_422),
.B(n_418),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_812),
.A2(n_844),
.B1(n_836),
.B2(n_828),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_829),
.A2(n_17),
.B(n_18),
.C(n_23),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_887),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_759),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_754),
.B(n_799),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_839),
.B(n_422),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_835),
.A2(n_422),
.B1(n_418),
.B2(n_416),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_778),
.B(n_856),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_802),
.A2(n_418),
.B(n_416),
.C(n_27),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_843),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_784),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_813),
.A2(n_418),
.B(n_416),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_839),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_821),
.B(n_418),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_771),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_800),
.A2(n_418),
.B(n_416),
.C(n_28),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_SL g962 ( 
.A1(n_730),
.A2(n_69),
.B(n_136),
.C(n_134),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_762),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_811),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_728),
.B(n_23),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_743),
.B(n_416),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_728),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_762),
.B(n_87),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_877),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_816),
.A2(n_416),
.B(n_88),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_747),
.A2(n_416),
.B1(n_39),
.B2(n_41),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_744),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_811),
.B(n_91),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_753),
.A2(n_75),
.B(n_117),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_784),
.Y(n_975)
);

OA22x2_ASAP7_75t_L g976 ( 
.A1(n_773),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_760),
.B(n_47),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_724),
.A2(n_68),
.B(n_111),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_787),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_790),
.B(n_101),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_775),
.A2(n_60),
.B(n_110),
.Y(n_981)
);

BUFx6f_ASAP7_75t_SL g982 ( 
.A(n_773),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_773),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_SL g984 ( 
.A1(n_779),
.A2(n_127),
.B(n_107),
.C(n_106),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_820),
.B(n_103),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_811),
.B(n_751),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_838),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_L g988 ( 
.A1(n_830),
.A2(n_56),
.B(n_59),
.C(n_729),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_724),
.A2(n_726),
.B(n_727),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_752),
.A2(n_727),
.B(n_726),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_764),
.B(n_755),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_SL g992 ( 
.A1(n_863),
.A2(n_874),
.B(n_867),
.C(n_853),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_851),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_765),
.A2(n_767),
.B(n_881),
.Y(n_994)
);

AO32x2_ASAP7_75t_L g995 ( 
.A1(n_777),
.A2(n_781),
.A3(n_806),
.B1(n_825),
.B2(n_822),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_881),
.A2(n_756),
.B(n_870),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_866),
.B(n_859),
.C(n_876),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_847),
.B(n_758),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_763),
.B(n_811),
.Y(n_999)
);

OR2x6_ASAP7_75t_L g1000 ( 
.A(n_851),
.B(n_735),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_811),
.B(n_837),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_792),
.Y(n_1002)
);

AO32x1_ASAP7_75t_L g1003 ( 
.A1(n_882),
.A2(n_841),
.A3(n_798),
.B1(n_793),
.B2(n_817),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_731),
.B(n_878),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_735),
.A2(n_826),
.B(n_833),
.Y(n_1005)
);

AO21x2_ASAP7_75t_L g1006 ( 
.A1(n_772),
.A2(n_840),
.B(n_886),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_824),
.A2(n_804),
.B(n_884),
.C(n_885),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_801),
.B(n_886),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_885),
.A2(n_888),
.B(n_872),
.C(n_871),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_898),
.A2(n_888),
.B(n_871),
.C(n_869),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_898),
.B(n_869),
.Y(n_1011)
);

AOI221xp5_ASAP7_75t_SL g1012 ( 
.A1(n_890),
.A2(n_858),
.B1(n_861),
.B2(n_862),
.C(n_846),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_932),
.A2(n_795),
.B(n_803),
.Y(n_1013)
);

AO32x2_ASAP7_75t_L g1014 ( 
.A1(n_971),
.A2(n_857),
.A3(n_850),
.B1(n_848),
.B2(n_846),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_902),
.A2(n_794),
.B(n_865),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_990),
.A2(n_848),
.B(n_850),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_988),
.A2(n_873),
.B(n_854),
.C(n_849),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_927),
.B(n_769),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1004),
.A2(n_845),
.B(n_815),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_893),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_946),
.A2(n_818),
.B(n_823),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_996),
.A2(n_805),
.B(n_807),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_994),
.A2(n_810),
.B(n_1005),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_953),
.A2(n_985),
.B1(n_891),
.B2(n_998),
.Y(n_1024)
);

AO31x2_ASAP7_75t_L g1025 ( 
.A1(n_934),
.A2(n_961),
.A3(n_946),
.B(n_954),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_926),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_935),
.A2(n_925),
.B(n_989),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_950),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_931),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_967),
.B(n_921),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_960),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_942),
.A2(n_1008),
.B(n_1000),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_897),
.A2(n_979),
.B1(n_907),
.B2(n_911),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_895),
.A2(n_1009),
.B(n_981),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_914),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_962),
.A2(n_984),
.B(n_973),
.C(n_977),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_906),
.A2(n_971),
.A3(n_1002),
.B(n_903),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_924),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_958),
.B(n_901),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_889),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_945),
.A2(n_957),
.B(n_938),
.Y(n_1041)
);

AO31x2_ASAP7_75t_L g1042 ( 
.A1(n_903),
.A2(n_952),
.A3(n_970),
.B(n_986),
.Y(n_1042)
);

OAI22x1_ASAP7_75t_L g1043 ( 
.A1(n_965),
.A2(n_985),
.B1(n_983),
.B2(n_913),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_997),
.A2(n_1007),
.B(n_910),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_916),
.A2(n_937),
.B(n_972),
.C(n_947),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_975),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_899),
.B(n_991),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_909),
.B(n_912),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_900),
.A2(n_987),
.B(n_997),
.C(n_941),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_899),
.B(n_991),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_936),
.B(n_1001),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1000),
.A2(n_966),
.B(n_944),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_939),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_978),
.A2(n_952),
.B(n_964),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_972),
.A2(n_922),
.B(n_951),
.C(n_920),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1000),
.A2(n_944),
.B(n_1006),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_974),
.A2(n_948),
.B(n_930),
.C(n_956),
.Y(n_1058)
);

AO31x2_ASAP7_75t_L g1059 ( 
.A1(n_1003),
.A2(n_896),
.A3(n_975),
.B(n_1006),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_956),
.B(n_949),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_904),
.A2(n_968),
.B(n_915),
.C(n_918),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_894),
.B(n_905),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1003),
.A2(n_949),
.B(n_905),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_963),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_915),
.B(n_955),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_933),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_923),
.A2(n_976),
.B1(n_943),
.B2(n_982),
.Y(n_1067)
);

AOI221x1_ASAP7_75t_L g1068 ( 
.A1(n_995),
.A2(n_931),
.B1(n_940),
.B2(n_943),
.C(n_959),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_917),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_969),
.B(n_928),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_959),
.B(n_931),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_919),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_999),
.A2(n_940),
.B(n_963),
.Y(n_1073)
);

AOI21x1_ASAP7_75t_L g1074 ( 
.A1(n_995),
.A2(n_959),
.B(n_980),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_993),
.A2(n_940),
.B(n_995),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_980),
.A2(n_963),
.B(n_982),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_990),
.A2(n_841),
.B(n_996),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_898),
.B(n_597),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_992),
.A2(n_814),
.B(n_785),
.C(n_647),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_785),
.B1(n_898),
.B2(n_814),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_898),
.B(n_785),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_992),
.A2(n_814),
.B(n_785),
.C(n_647),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_971),
.A2(n_990),
.B1(n_785),
.B2(n_814),
.C(n_954),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_937),
.A2(n_814),
.B1(n_646),
.B2(n_785),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_893),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_893),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_950),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_992),
.A2(n_932),
.B(n_716),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_992),
.A2(n_932),
.B(n_716),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_898),
.B(n_785),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_893),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_992),
.A2(n_785),
.B(n_892),
.C(n_962),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_927),
.B(n_929),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_967),
.B(n_921),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_990),
.A2(n_841),
.B(n_996),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_992),
.A2(n_932),
.B(n_716),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_992),
.A2(n_814),
.B(n_785),
.C(n_647),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_890),
.A2(n_785),
.B1(n_898),
.B2(n_814),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_927),
.B(n_929),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_932),
.A2(n_946),
.B(n_997),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_898),
.B(n_785),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_898),
.B(n_597),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_932),
.A2(n_946),
.B(n_997),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_960),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_990),
.A2(n_841),
.B(n_996),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_937),
.B(n_814),
.C(n_785),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_958),
.B(n_619),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_990),
.A2(n_841),
.B(n_996),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_990),
.A2(n_989),
.B(n_996),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_932),
.A2(n_946),
.B(n_997),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_898),
.A2(n_814),
.B(n_785),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_898),
.B(n_785),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_898),
.B(n_785),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_963),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_898),
.B(n_785),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_990),
.A2(n_841),
.B(n_996),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_927),
.B(n_929),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_992),
.A2(n_932),
.B(n_716),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_890),
.A2(n_785),
.B1(n_898),
.B2(n_814),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_898),
.A2(n_785),
.B(n_814),
.C(n_597),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_958),
.B(n_619),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_SL g1122 ( 
.A(n_937),
.B(n_785),
.C(n_814),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_SL g1123 ( 
.A(n_908),
.B(n_960),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_898),
.A2(n_785),
.B(n_814),
.C(n_597),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_953),
.A2(n_814),
.B1(n_785),
.B2(n_319),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_927),
.B(n_929),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_992),
.A2(n_932),
.B(n_716),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_L g1128 ( 
.A(n_975),
.B(n_956),
.Y(n_1128)
);

BUFx8_ASAP7_75t_L g1129 ( 
.A(n_982),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1106),
.A2(n_1119),
.B1(n_1098),
.B2(n_1080),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_1031),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1080),
.A2(n_1119),
.B1(n_1098),
.B2(n_1065),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1122),
.A2(n_1084),
.B1(n_1111),
.B2(n_1125),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1093),
.A2(n_1117),
.B(n_1099),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1026),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1024),
.A2(n_1081),
.B1(n_1101),
.B2(n_1113),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1029),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_1104),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1112),
.A2(n_1115),
.B1(n_1090),
.B2(n_1044),
.Y(n_1139)
);

CKINVDCx11_ASAP7_75t_R g1140 ( 
.A(n_1040),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1078),
.B(n_1102),
.Y(n_1141)
);

INVx6_ASAP7_75t_L g1142 ( 
.A(n_1029),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1072),
.Y(n_1143)
);

INVx6_ASAP7_75t_L g1144 ( 
.A(n_1029),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1044),
.A2(n_1110),
.B1(n_1103),
.B2(n_1100),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1045),
.A2(n_1120),
.B(n_1124),
.Y(n_1146)
);

CKINVDCx11_ASAP7_75t_R g1147 ( 
.A(n_1028),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1093),
.B(n_1099),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1129),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1117),
.B(n_1126),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1129),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1100),
.A2(n_1103),
.B1(n_1110),
.B2(n_1043),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1107),
.B(n_1121),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1079),
.A2(n_1097),
.B(n_1082),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_SL g1156 ( 
.A(n_1055),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1028),
.Y(n_1157)
);

INVx5_ASAP7_75t_SL g1158 ( 
.A(n_1030),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1083),
.A2(n_1050),
.B1(n_1047),
.B2(n_1068),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1033),
.A2(n_1011),
.B1(n_1050),
.B2(n_1047),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1069),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1085),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1046),
.B(n_1076),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_SL g1164 ( 
.A(n_1030),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_1094),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1033),
.A2(n_1067),
.B1(n_1018),
.B2(n_1051),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1038),
.A2(n_1053),
.B1(n_1091),
.B2(n_1086),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1087),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1039),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1048),
.Y(n_1170)
);

CKINVDCx11_ASAP7_75t_R g1171 ( 
.A(n_1114),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1064),
.Y(n_1172)
);

INVx6_ASAP7_75t_L g1173 ( 
.A(n_1123),
.Y(n_1173)
);

INVx6_ASAP7_75t_L g1174 ( 
.A(n_1064),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1071),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1062),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1075),
.A2(n_1057),
.B1(n_1052),
.B2(n_1066),
.Y(n_1177)
);

CKINVDCx12_ASAP7_75t_R g1178 ( 
.A(n_1073),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1074),
.A2(n_1071),
.B1(n_1046),
.B2(n_1128),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1032),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1014),
.Y(n_1181)
);

INVx6_ASAP7_75t_L g1182 ( 
.A(n_1058),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1014),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1010),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1021),
.A2(n_1127),
.B1(n_1118),
.B2(n_1088),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1021),
.A2(n_1096),
.B1(n_1089),
.B2(n_1019),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1037),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_1060),
.B1(n_1063),
.B2(n_1016),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1059),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1041),
.A2(n_1013),
.B1(n_1054),
.B2(n_1027),
.Y(n_1190)
);

BUFx8_ASAP7_75t_SL g1191 ( 
.A(n_1109),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1015),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1092),
.Y(n_1193)
);

INVx6_ASAP7_75t_L g1194 ( 
.A(n_1012),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_1023),
.B1(n_1061),
.B2(n_1116),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1022),
.Y(n_1196)
);

BUFx4_ASAP7_75t_SL g1197 ( 
.A(n_1012),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1036),
.A2(n_1056),
.B1(n_1025),
.B2(n_1017),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1059),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1025),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1042),
.B(n_1077),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1042),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1042),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1095),
.Y(n_1204)
);

AOI22x1_ASAP7_75t_SL g1205 ( 
.A1(n_1105),
.A2(n_919),
.B1(n_401),
.B2(n_590),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1108),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1029),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1026),
.Y(n_1208)
);

BUFx8_ASAP7_75t_L g1209 ( 
.A(n_1031),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1031),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1125),
.A2(n_785),
.B1(n_1106),
.B2(n_1024),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1122),
.A2(n_814),
.B1(n_1106),
.B2(n_785),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1122),
.A2(n_814),
.B1(n_1106),
.B2(n_785),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1026),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1125),
.A2(n_785),
.B1(n_1106),
.B2(n_1024),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1081),
.B(n_1090),
.Y(n_1217)
);

INVx6_ASAP7_75t_L g1218 ( 
.A(n_1029),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1106),
.A2(n_814),
.B1(n_646),
.B2(n_785),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1031),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1026),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1122),
.A2(n_814),
.B1(n_1106),
.B2(n_785),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1020),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1026),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1078),
.B(n_1102),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1122),
.A2(n_814),
.B1(n_1106),
.B2(n_785),
.Y(n_1226)
);

BUFx8_ASAP7_75t_SL g1227 ( 
.A(n_1031),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1029),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_SL g1229 ( 
.A(n_1070),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1122),
.A2(n_814),
.B1(n_1106),
.B2(n_785),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1125),
.A2(n_785),
.B1(n_1106),
.B2(n_1024),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_1125),
.B1(n_814),
.B2(n_785),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1125),
.A2(n_785),
.B1(n_1106),
.B2(n_1024),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1125),
.A2(n_814),
.B(n_1084),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1081),
.B(n_1090),
.Y(n_1235)
);

INVx6_ASAP7_75t_L g1236 ( 
.A(n_1029),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1029),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1020),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1187),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1133),
.A2(n_1219),
.B1(n_1234),
.B2(n_1232),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1175),
.B(n_1151),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1151),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1195),
.A2(n_1190),
.B(n_1185),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1132),
.B(n_1153),
.Y(n_1245)
);

BUFx2_ASAP7_75t_SL g1246 ( 
.A(n_1164),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1169),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1155),
.A2(n_1201),
.B(n_1198),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1203),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1180),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1135),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1141),
.B(n_1225),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1223),
.Y(n_1253)
);

OR2x2_ASAP7_75t_SL g1254 ( 
.A(n_1173),
.B(n_1194),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1154),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1211),
.A2(n_1231),
.B1(n_1233),
.B2(n_1216),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1146),
.B(n_1136),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_1173),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1153),
.B(n_1145),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1202),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1145),
.B(n_1130),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1200),
.B(n_1160),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1183),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1183),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1175),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1175),
.B(n_1238),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1217),
.B(n_1235),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1194),
.B(n_1238),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1140),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1184),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1170),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1176),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1166),
.B(n_1139),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1195),
.A2(n_1190),
.B(n_1185),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1166),
.B(n_1139),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1229),
.B(n_1208),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1162),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1214),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1226),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1165),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1186),
.A2(n_1206),
.B(n_1204),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1165),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1189),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_R g1284 ( 
.A(n_1138),
.B(n_1220),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1197),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1224),
.B(n_1136),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1186),
.A2(n_1206),
.B(n_1188),
.Y(n_1287)
);

AND2x2_ASAP7_75t_SL g1288 ( 
.A(n_1177),
.B(n_1133),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1147),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_R g1290 ( 
.A(n_1131),
.B(n_1210),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1134),
.Y(n_1291)
);

CKINVDCx6p67_ASAP7_75t_R g1292 ( 
.A(n_1152),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1199),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1163),
.B(n_1182),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1181),
.Y(n_1295)
);

BUFx4f_ASAP7_75t_SL g1296 ( 
.A(n_1157),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1159),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1212),
.A2(n_1230),
.B(n_1226),
.C(n_1222),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1159),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1182),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1177),
.B(n_1167),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1182),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1213),
.B(n_1192),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1196),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1179),
.A2(n_1221),
.B(n_1215),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1196),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1193),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1179),
.B(n_1158),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1191),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1178),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1173),
.A2(n_1172),
.B1(n_1164),
.B2(n_1135),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1291),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1243),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1241),
.A2(n_1161),
.B(n_1205),
.C(n_1168),
.Y(n_1314)
);

OAI21xp33_ASAP7_75t_L g1315 ( 
.A1(n_1256),
.A2(n_1149),
.B(n_1137),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1244),
.A2(n_1142),
.B(n_1236),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1255),
.B(n_1242),
.Y(n_1317)
);

INVx5_ASAP7_75t_SL g1318 ( 
.A(n_1292),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1257),
.B(n_1174),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1257),
.B(n_1171),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1309),
.A2(n_1156),
.B1(n_1237),
.B2(n_1144),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1258),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1242),
.B(n_1143),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1286),
.B(n_1142),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1288),
.A2(n_1144),
.B(n_1236),
.C(n_1207),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1308),
.B(n_1207),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1288),
.A2(n_1209),
.B1(n_1156),
.B2(n_1218),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1258),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1279),
.A2(n_1218),
.B1(n_1227),
.B2(n_1228),
.C(n_1298),
.Y(n_1329)
);

OR2x2_ASAP7_75t_SL g1330 ( 
.A(n_1309),
.B(n_1310),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1266),
.B(n_1262),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1288),
.A2(n_1245),
.B(n_1261),
.C(n_1291),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1277),
.B(n_1278),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1240),
.A2(n_1267),
.B(n_1248),
.Y(n_1335)
);

INVxp33_ASAP7_75t_L g1336 ( 
.A(n_1252),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1245),
.A2(n_1261),
.B(n_1275),
.C(n_1273),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1273),
.A2(n_1275),
.B(n_1259),
.C(n_1301),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_SL g1340 ( 
.A(n_1294),
.B(n_1308),
.Y(n_1340)
);

AOI211xp5_ASAP7_75t_L g1341 ( 
.A1(n_1297),
.A2(n_1299),
.B(n_1305),
.C(n_1310),
.Y(n_1341)
);

NOR2x1_ASAP7_75t_SL g1342 ( 
.A(n_1294),
.B(n_1248),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1247),
.B(n_1271),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_SL g1344 ( 
.A1(n_1300),
.A2(n_1302),
.B(n_1285),
.C(n_1307),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1244),
.A2(n_1274),
.B(n_1287),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1250),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1269),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1248),
.A2(n_1294),
.B(n_1300),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1272),
.B(n_1303),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1265),
.B(n_1301),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1274),
.A2(n_1281),
.B(n_1287),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1285),
.A2(n_1246),
.B1(n_1297),
.B2(n_1299),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1254),
.A2(n_1303),
.B1(n_1307),
.B2(n_1302),
.Y(n_1353)
);

AOI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1270),
.A2(n_1268),
.B1(n_1311),
.B2(n_1283),
.C(n_1246),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1312),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1345),
.B(n_1295),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1313),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1335),
.B(n_1270),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1313),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1351),
.B(n_1249),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1334),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1316),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1334),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1316),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1346),
.B(n_1283),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1342),
.B(n_1239),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1336),
.B(n_1254),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1333),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_L g1370 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1349),
.B(n_1250),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1339),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1339),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1320),
.A2(n_1353),
.B1(n_1332),
.B2(n_1318),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1343),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1325),
.B(n_1253),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1350),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1358),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1377),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1356),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1359),
.B(n_1355),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1359),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1361),
.A2(n_1293),
.B(n_1260),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1375),
.A2(n_1329),
.B1(n_1315),
.B2(n_1320),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1368),
.B(n_1336),
.Y(n_1387)
);

AOI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1375),
.A2(n_1341),
.B(n_1314),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1356),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1356),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1377),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1360),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1372),
.B(n_1340),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1369),
.B(n_1338),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1372),
.B(n_1331),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1368),
.A2(n_1332),
.B1(n_1337),
.B2(n_1338),
.Y(n_1396)
);

NOR2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1377),
.B(n_1292),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1377),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1371),
.B(n_1366),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1370),
.B(n_1326),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1401)
);

OAI211xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1370),
.A2(n_1337),
.B(n_1354),
.C(n_1327),
.Y(n_1402)
);

AOI33xp33_ASAP7_75t_L g1403 ( 
.A1(n_1357),
.A2(n_1352),
.A3(n_1289),
.B1(n_1317),
.B2(n_1344),
.B3(n_1323),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1357),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1404),
.B(n_1363),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1381),
.B(n_1367),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1390),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1385),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1401),
.B(n_1363),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1385),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1391),
.B(n_1362),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1384),
.B(n_1363),
.Y(n_1412)
);

NAND4xp25_ASAP7_75t_L g1413 ( 
.A(n_1388),
.B(n_1386),
.C(n_1402),
.D(n_1396),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1384),
.B(n_1379),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1385),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1385),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1394),
.B(n_1379),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1388),
.A2(n_1344),
.B(n_1325),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1391),
.B(n_1364),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1391),
.B(n_1364),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1387),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1394),
.B(n_1376),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1391),
.B(n_1364),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1382),
.B(n_1365),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1382),
.B(n_1366),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1389),
.B(n_1366),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1398),
.B(n_1373),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1392),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1376),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1392),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1390),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1380),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1398),
.B(n_1373),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1430),
.B(n_1383),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1406),
.B(n_1398),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1413),
.B(n_1284),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1429),
.Y(n_1438)
);

AOI21xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1413),
.A2(n_1396),
.B(n_1269),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1429),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1411),
.B(n_1398),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1423),
.B(n_1389),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1419),
.A2(n_1402),
.B(n_1386),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1411),
.B(n_1381),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1423),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1422),
.A2(n_1400),
.B1(n_1381),
.B2(n_1347),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1429),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1411),
.B(n_1381),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1431),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1407),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1431),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1420),
.B(n_1381),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1418),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1430),
.B(n_1383),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1431),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1418),
.B(n_1347),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

NOR3xp33_ASAP7_75t_L g1458 ( 
.A(n_1419),
.B(n_1387),
.C(n_1403),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1407),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1420),
.B(n_1393),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1414),
.B(n_1383),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1420),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1414),
.B(n_1399),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1432),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1426),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1421),
.B(n_1393),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1432),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1412),
.B(n_1399),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1405),
.A2(n_1378),
.B(n_1319),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1426),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1421),
.B(n_1393),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1424),
.B(n_1397),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1424),
.B(n_1397),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1474),
.B(n_1428),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1443),
.B(n_1428),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1467),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1456),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1458),
.B(n_1434),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1467),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1474),
.B(n_1434),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1453),
.B(n_1403),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1438),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1436),
.B(n_1406),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1475),
.B(n_1406),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1475),
.B(n_1409),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1440),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1450),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1439),
.B(n_1369),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1462),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1441),
.B(n_1409),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1440),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1497)
);

NOR2x1_ASAP7_75t_L g1498 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1395),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1444),
.B(n_1409),
.Y(n_1500)
);

OAI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1446),
.A2(n_1400),
.B1(n_1412),
.B2(n_1425),
.C(n_1371),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1447),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1448),
.B(n_1409),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1442),
.B(n_1395),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1459),
.B(n_1405),
.C(n_1319),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1435),
.B(n_1290),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1446),
.A2(n_1400),
.B1(n_1378),
.B2(n_1318),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1447),
.Y(n_1509)
);

NAND2x1_ASAP7_75t_L g1510 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1435),
.B(n_1427),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1492),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1498),
.A2(n_1464),
.B(n_1436),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1498),
.Y(n_1514)
);

AOI31xp33_ASAP7_75t_L g1515 ( 
.A1(n_1494),
.A2(n_1448),
.A3(n_1452),
.B(n_1276),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_1479),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1484),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1492),
.B(n_1436),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1497),
.Y(n_1519)
);

OAI211xp5_ASAP7_75t_L g1520 ( 
.A1(n_1481),
.A2(n_1468),
.B(n_1452),
.C(n_1461),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1486),
.A2(n_1400),
.B1(n_1454),
.B2(n_1461),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1479),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1487),
.Y(n_1525)
);

AOI222xp33_ASAP7_75t_L g1526 ( 
.A1(n_1506),
.A2(n_1405),
.B1(n_1442),
.B2(n_1476),
.C1(n_1470),
.C2(n_1468),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1497),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1482),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1476),
.Y(n_1529)
);

AOI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1507),
.A2(n_1454),
.B(n_1472),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1493),
.B(n_1460),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1482),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1477),
.B(n_1460),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1501),
.B(n_1296),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1506),
.A2(n_1321),
.B1(n_1400),
.B2(n_1324),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1508),
.A2(n_1463),
.B(n_1472),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1514),
.A2(n_1508),
.B(n_1482),
.Y(n_1537)
);

AOI21xp33_ASAP7_75t_L g1538 ( 
.A1(n_1513),
.A2(n_1485),
.B(n_1510),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_L g1539 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1485),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1512),
.B(n_1477),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1516),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1483),
.Y(n_1544)
);

INVxp33_ASAP7_75t_L g1545 ( 
.A(n_1531),
.Y(n_1545)
);

INVxp33_ASAP7_75t_L g1546 ( 
.A(n_1534),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1518),
.Y(n_1547)
);

OAI21xp33_ASAP7_75t_L g1548 ( 
.A1(n_1529),
.A2(n_1499),
.B(n_1483),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1511),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1530),
.B(n_1502),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1526),
.A2(n_1490),
.B1(n_1495),
.B2(n_1489),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

OAI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1536),
.A2(n_1490),
.B(n_1489),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1536),
.A2(n_1510),
.B(n_1488),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1524),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1543),
.B(n_1524),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1549),
.A2(n_1520),
.B1(n_1518),
.B2(n_1533),
.Y(n_1558)
);

XNOR2x1_ASAP7_75t_L g1559 ( 
.A(n_1539),
.B(n_1535),
.Y(n_1559)
);

XNOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1540),
.B(n_1521),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1545),
.B(n_1533),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1546),
.A2(n_1400),
.B1(n_1511),
.B2(n_1532),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1537),
.A2(n_1532),
.B(n_1528),
.C(n_1525),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1544),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1544),
.B(n_1495),
.Y(n_1565)
);

NOR2x1p5_ASAP7_75t_SL g1566 ( 
.A(n_1555),
.B(n_1528),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1558),
.A2(n_1551),
.B1(n_1552),
.B2(n_1547),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1569)
);

NOR3x1_ASAP7_75t_L g1570 ( 
.A(n_1563),
.B(n_1537),
.C(n_1550),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1559),
.B(n_1557),
.C(n_1563),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1560),
.A2(n_1554),
.B(n_1538),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1561),
.B(n_1553),
.C(n_1565),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1566),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1562),
.B(n_1523),
.C(n_1517),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1564),
.B(n_1517),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1571),
.B(n_1523),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1567),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1568),
.A2(n_1488),
.B1(n_1525),
.B2(n_1491),
.Y(n_1579)
);

AOI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1572),
.A2(n_1509),
.B1(n_1487),
.B2(n_1491),
.C(n_1503),
.Y(n_1580)
);

AOI211xp5_ASAP7_75t_L g1581 ( 
.A1(n_1574),
.A2(n_1488),
.B(n_1509),
.C(n_1496),
.Y(n_1581)
);

AOI21xp33_ASAP7_75t_L g1582 ( 
.A1(n_1569),
.A2(n_1496),
.B(n_1503),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1575),
.A2(n_1488),
.B(n_1405),
.C(n_1500),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1579),
.A2(n_1573),
.B(n_1576),
.Y(n_1584)
);

AOI211xp5_ASAP7_75t_L g1585 ( 
.A1(n_1582),
.A2(n_1578),
.B(n_1581),
.C(n_1583),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1570),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1580),
.A2(n_1504),
.B1(n_1500),
.B2(n_1465),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1577),
.A2(n_1457),
.B(n_1471),
.C(n_1465),
.Y(n_1588)
);

NAND4xp25_ASAP7_75t_L g1589 ( 
.A(n_1579),
.B(n_1504),
.C(n_1505),
.D(n_1251),
.Y(n_1589)
);

OAI322xp33_ASAP7_75t_L g1590 ( 
.A1(n_1579),
.A2(n_1416),
.A3(n_1408),
.B1(n_1415),
.B2(n_1417),
.C1(n_1410),
.C2(n_1457),
.Y(n_1590)
);

NOR3xp33_ASAP7_75t_L g1591 ( 
.A(n_1584),
.B(n_1463),
.C(n_1471),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1586),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1585),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1588),
.Y(n_1594)
);

XOR2xp5_ASAP7_75t_L g1595 ( 
.A(n_1589),
.B(n_1318),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1592),
.A2(n_1591),
.B(n_1587),
.Y(n_1596)
);

AOI221x1_ASAP7_75t_L g1597 ( 
.A1(n_1593),
.A2(n_1594),
.B1(n_1595),
.B2(n_1590),
.C(n_1449),
.Y(n_1597)
);

OA22x2_ASAP7_75t_L g1598 ( 
.A1(n_1595),
.A2(n_1449),
.B1(n_1451),
.B2(n_1455),
.Y(n_1598)
);

OAI211xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1596),
.A2(n_1455),
.B(n_1451),
.C(n_1425),
.Y(n_1599)
);

OAI22x1_ASAP7_75t_L g1600 ( 
.A1(n_1599),
.A2(n_1597),
.B1(n_1598),
.B2(n_1473),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1600),
.Y(n_1601)
);

OAI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1600),
.A2(n_1473),
.B(n_1466),
.Y(n_1602)
);

AOI22x1_ASAP7_75t_L g1603 ( 
.A1(n_1601),
.A2(n_1282),
.B1(n_1280),
.B2(n_1466),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1602),
.A2(n_1425),
.B1(n_1427),
.B2(n_1433),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1603),
.B(n_1604),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1603),
.B(n_1433),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1605),
.A2(n_1408),
.B1(n_1410),
.B2(n_1417),
.Y(n_1607)
);

OAI321xp33_ASAP7_75t_L g1608 ( 
.A1(n_1607),
.A2(n_1606),
.A3(n_1408),
.B1(n_1415),
.B2(n_1417),
.C(n_1416),
.Y(n_1608)
);

BUFx4_ASAP7_75t_R g1609 ( 
.A(n_1608),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_R g1610 ( 
.A1(n_1609),
.A2(n_1258),
.B1(n_1410),
.B2(n_1415),
.C(n_1417),
.Y(n_1610)
);

AOI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1610),
.A2(n_1328),
.B(n_1322),
.C(n_1282),
.Y(n_1611)
);


endmodule