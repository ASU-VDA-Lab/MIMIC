module fake_jpeg_13326_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_8),
.B(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_45),
.B1(n_38),
.B2(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_12),
.B1(n_25),
.B2(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_34),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.C(n_38),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_70),
.B1(n_72),
.B2(n_13),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_3),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_9),
.C(n_10),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_56),
.B1(n_60),
.B2(n_48),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_74),
.B1(n_8),
.B2(n_9),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_81),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_11),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_68),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_76),
.B1(n_65),
.B2(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_70),
.B1(n_87),
.B2(n_89),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_92),
.B(n_86),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_94),
.Y(n_95)
);

AOI31xp67_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_78),
.A3(n_86),
.B(n_21),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_96),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_18),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_20),
.Y(n_99)
);


endmodule