module fake_jpeg_21724_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_21),
.B1(n_29),
.B2(n_34),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_29),
.B1(n_35),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_35),
.B1(n_24),
.B2(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_33),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_71),
.Y(n_115)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_30),
.C(n_32),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_30),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_45),
.C(n_38),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_109),
.C(n_31),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_67),
.A3(n_62),
.B1(n_53),
.B2(n_63),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_32),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_36),
.B1(n_39),
.B2(n_45),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_36),
.B1(n_37),
.B2(n_17),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_37),
.B1(n_36),
.B2(n_17),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_92),
.B1(n_96),
.B2(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_30),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_40),
.B1(n_23),
.B2(n_27),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_102),
.Y(n_134)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_33),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_15),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_48),
.B(n_33),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_31),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_40),
.B(n_32),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_27),
.Y(n_135)
);

BUFx2_ASAP7_75t_SL g108 ( 
.A(n_49),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_31),
.C(n_27),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_113),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_124),
.B1(n_130),
.B2(n_105),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_31),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_105),
.B1(n_70),
.B2(n_80),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_32),
.B(n_30),
.Y(n_122)
);

OR2x4_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_125),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_68),
.B1(n_92),
.B2(n_86),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_R g153 ( 
.A(n_125),
.B(n_137),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_40),
.B1(n_27),
.B2(n_26),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_25),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_10),
.Y(n_169)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_159),
.C(n_110),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_91),
.B1(n_86),
.B2(n_96),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_150),
.B1(n_162),
.B2(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_79),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_81),
.B1(n_85),
.B2(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_165),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_81),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_157),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_119),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_98),
.C(n_88),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_93),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_164),
.Y(n_202)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_74),
.B1(n_26),
.B2(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_100),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_26),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_113),
.B(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_25),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_123),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_186),
.B1(n_145),
.B2(n_163),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_164),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_180),
.A2(n_181),
.B1(n_126),
.B2(n_161),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_133),
.B1(n_125),
.B2(n_110),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_125),
.B(n_123),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_191),
.B(n_166),
.Y(n_220)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_115),
.B1(n_138),
.B2(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_137),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_11),
.C(n_16),
.Y(n_227)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_203),
.C(n_126),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_137),
.C(n_131),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_157),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_212),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_144),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_217),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_146),
.B1(n_149),
.B2(n_167),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_230),
.B1(n_191),
.B2(n_199),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_202),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_221),
.A2(n_223),
.B(n_231),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_136),
.B(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_159),
.B(n_147),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_203),
.C(n_176),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

OA21x2_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_196),
.B(n_8),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_200),
.B1(n_195),
.B2(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_133),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_25),
.B(n_8),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_239),
.B1(n_243),
.B2(n_205),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_209),
.B1(n_210),
.B2(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_249),
.C(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_215),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_253),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_194),
.B1(n_202),
.B2(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_230),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_194),
.B(n_179),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_251),
.B(n_219),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_197),
.C(n_196),
.Y(n_249)
);

NOR4xp25_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_185),
.C(n_183),
.D(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_225),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_220),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_217),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_263),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_218),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_231),
.B1(n_209),
.B2(n_210),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_232),
.B1(n_244),
.B2(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_229),
.C(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.C(n_271),
.Y(n_281)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_222),
.C(n_221),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_222),
.C(n_205),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_235),
.B1(n_248),
.B2(n_233),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_0),
.B(n_1),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_282),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_267),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_268),
.CI(n_254),
.CON(n_285),
.SN(n_285)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_234),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_240),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_284),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_269),
.B(n_274),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_283),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_261),
.B1(n_260),
.B2(n_236),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_273),
.B1(n_285),
.B2(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_264),
.C(n_185),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_298),
.C(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_0),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_11),
.C(n_15),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_303),
.B(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_279),
.C(n_276),
.Y(n_303)
);

AOI221xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.C(n_12),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_292),
.Y(n_305)
);

NAND4xp25_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_291),
.C(n_293),
.D(n_295),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_301),
.B(n_303),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_288),
.B(n_298),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_310),
.B(n_312),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_297),
.B(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_311),
.B(n_5),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_4),
.B(n_5),
.Y(n_315)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_7),
.B(n_12),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_7),
.B1(n_13),
.B2(n_16),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_13),
.Y(n_321)
);


endmodule