module fake_netlist_1_713_n_41 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
BUFx8_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_9), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_13), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_1), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_19), .B(n_0), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_16), .Y(n_26) );
AOI221xp5_ASAP7_75t_SL g27 ( .A1(n_18), .A2(n_21), .B1(n_20), .B2(n_17), .C(n_22), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_23), .Y(n_28) );
O2A1O1Ixp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_17), .B(n_22), .C(n_16), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_6), .B(n_14), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_26), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_24), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_24), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_33), .B(n_24), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_15), .B1(n_30), .B2(n_25), .C1(n_26), .C2(n_31), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_15), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NAND4xp25_ASAP7_75t_L g38 ( .A(n_36), .B(n_2), .C(n_4), .D(n_5), .Y(n_38) );
OR2x2_ASAP7_75t_L g39 ( .A(n_38), .B(n_37), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
endmodule