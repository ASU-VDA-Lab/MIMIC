module fake_netlist_1_12595_n_701 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_701);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_701;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_17), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_18), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_53), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_26), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_80), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_59), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_73), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_44), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_64), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_57), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_81), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_84), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_24), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_49), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_25), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_95), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_55), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_93), .B(n_3), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_5), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_28), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_97), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_90), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_43), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_31), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_14), .Y(n_131) );
BUFx8_ASAP7_75t_SL g132 ( .A(n_2), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_1), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_6), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_58), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_48), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_46), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_88), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_91), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_3), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_34), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_50), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_5), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_52), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_15), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g148 ( .A1(n_103), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_105), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_105), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_133), .B(n_0), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_105), .Y(n_154) );
NOR2x1_ASAP7_75t_L g155 ( .A(n_114), .B(n_21), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_106), .B(n_4), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_106), .B(n_4), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_105), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_147), .B(n_117), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_157), .B(n_113), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_160), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_160), .B(n_119), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_147), .B(n_118), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_152), .A2(n_125), .B1(n_124), .B2(n_143), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_152), .B(n_120), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_158), .B(n_121), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_163), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_153), .B(n_129), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_161), .B(n_145), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_159), .B(n_135), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_166), .B(n_153), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_183), .B(n_111), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_177), .B(n_111), .Y(n_197) );
NAND2x1_ASAP7_75t_L g198 ( .A(n_181), .B(n_137), .Y(n_198) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_183), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_174), .B(n_155), .C(n_141), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_184), .A2(n_140), .B1(n_148), .B2(n_145), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_188), .B(n_136), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_188), .B(n_136), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_169), .B(n_138), .Y(n_206) );
BUFx8_ASAP7_75t_L g207 ( .A(n_168), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_168), .B(n_138), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_167), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_175), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g212 ( .A(n_174), .B(n_144), .C(n_102), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_184), .A2(n_139), .B1(n_109), .B2(n_110), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_139), .B1(n_109), .B2(n_110), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_169), .B(n_142), .Y(n_215) );
NAND3xp33_ASAP7_75t_SL g216 ( .A(n_187), .B(n_126), .C(n_142), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_184), .B(n_116), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_187), .B(n_128), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_187), .B(n_122), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_169), .B(n_127), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_184), .B(n_130), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_184), .B(n_108), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_184), .B(n_126), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_184), .B(n_123), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_194), .B(n_175), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_203), .B(n_184), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_173), .B(n_176), .C(n_165), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_223), .A2(n_173), .B1(n_176), .B2(n_165), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_205), .B(n_169), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_196), .B(n_169), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_208), .B(n_179), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_179), .B(n_180), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_218), .B(n_132), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_200), .B(n_180), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_213), .A2(n_108), .B1(n_149), .B2(n_150), .Y(n_239) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_198), .A2(n_195), .B(n_206), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_222), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_199), .B(n_108), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_219), .B(n_6), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_182), .B(n_172), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g246 ( .A(n_207), .B(n_108), .C(n_190), .Y(n_246) );
INVx5_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_191), .Y(n_248) );
OAI321xp33_ASAP7_75t_L g249 ( .A1(n_201), .A2(n_149), .A3(n_150), .B1(n_154), .B2(n_162), .C(n_108), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_216), .A2(n_149), .B1(n_150), .B2(n_154), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_215), .A2(n_190), .B(n_185), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_209), .B(n_7), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_201), .B(n_192), .C(n_212), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_225), .A2(n_214), .B1(n_212), .B2(n_209), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_254), .Y(n_258) );
AO31x2_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_224), .A3(n_204), .B(n_211), .Y(n_259) );
AOI21xp33_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_207), .B(n_197), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_220), .B(n_221), .Y(n_261) );
BUFx4f_ASAP7_75t_SL g262 ( .A(n_254), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_207), .B1(n_217), .B2(n_202), .Y(n_264) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_234), .A2(n_211), .A3(n_204), .B(n_185), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_237), .A2(n_172), .B(n_182), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_236), .A2(n_222), .B1(n_149), .B2(n_150), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_226), .A2(n_172), .B(n_182), .Y(n_268) );
OAI21x1_ASAP7_75t_SL g269 ( .A1(n_251), .A2(n_222), .B(n_8), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_233), .B(n_243), .C(n_239), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_178), .B(n_170), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_178), .B(n_170), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_229), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
AO31x2_ASAP7_75t_L g275 ( .A1(n_235), .A2(n_170), .A3(n_178), .B(n_162), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_238), .B(n_7), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_250), .B(n_8), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_251), .B(n_150), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_244), .A2(n_186), .B(n_189), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_279), .A2(n_249), .B(n_242), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_274), .B(n_263), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_279), .A2(n_270), .B(n_256), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_273), .B(n_238), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_276), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
BUFx8_ASAP7_75t_SL g286 ( .A(n_277), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_271), .A2(n_240), .B(n_253), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_246), .B(n_252), .Y(n_288) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_269), .A2(n_255), .B(n_248), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_268), .A2(n_241), .B(n_162), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_278), .A2(n_186), .B(n_189), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_258), .A2(n_241), .B(n_245), .C(n_247), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_264), .A2(n_154), .B(n_251), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_259), .B(n_232), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_257), .A2(n_154), .B(n_247), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_265), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_259), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_260), .A2(n_245), .B(n_247), .C(n_232), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_285), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_295), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
OA21x2_ASAP7_75t_L g304 ( .A1(n_282), .A2(n_272), .B(n_266), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_285), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_275), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_286), .A2(n_262), .B1(n_267), .B2(n_278), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
OAI21xp5_ASAP7_75t_L g311 ( .A1(n_282), .A2(n_247), .B(n_189), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_298), .A2(n_275), .B(n_154), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_298), .A2(n_275), .B(n_247), .Y(n_313) );
AO21x1_ASAP7_75t_SL g314 ( .A1(n_297), .A2(n_232), .B(n_61), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_297), .B(n_9), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_283), .B(n_232), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_9), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_294), .B(n_60), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_295), .A2(n_284), .B(n_299), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_298), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_283), .B(n_10), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_299), .B(n_10), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_296), .A2(n_11), .B(n_12), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_294), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_302), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_303), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_316), .B(n_284), .C(n_281), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_327), .B(n_294), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_327), .B(n_296), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_327), .B(n_289), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_309), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_307), .B(n_296), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_316), .B(n_290), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_322), .B(n_286), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_307), .B(n_296), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_309), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_307), .B(n_296), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_310), .B(n_293), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_305), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_321), .B(n_293), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_293), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_322), .B(n_289), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_321), .B(n_293), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_320), .B(n_289), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_306), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_320), .A2(n_287), .B(n_300), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_309), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_325), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_325), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_333), .B(n_309), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_329), .B(n_324), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_338), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_329), .B(n_324), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_333), .B(n_312), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_336), .B(n_312), .Y(n_381) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_332), .B(n_326), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_340), .B(n_312), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_340), .B(n_312), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_340), .B(n_312), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_343), .B(n_281), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_336), .B(n_319), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_347), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_352), .B(n_324), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_330), .Y(n_396) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_332), .B(n_323), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_344), .B(n_326), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_354), .B(n_318), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_344), .B(n_326), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_344), .B(n_326), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_355), .B(n_318), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_349), .B(n_326), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_328), .Y(n_405) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_342), .B(n_319), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_349), .B(n_319), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_349), .B(n_319), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_328), .B(n_319), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_331), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_334), .B(n_319), .Y(n_414) );
BUFx2_ASAP7_75t_SL g415 ( .A(n_339), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_334), .B(n_313), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_334), .B(n_313), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_331), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_356), .B(n_313), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_371), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_342), .B(n_308), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_335), .B(n_313), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_356), .B(n_313), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_335), .B(n_317), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_356), .B(n_317), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_358), .B(n_317), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_358), .B(n_293), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_365), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_339), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_429), .B(n_365), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_413), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_429), .B(n_365), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_430), .B(n_342), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_393), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_383), .B(n_358), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_375), .B(n_335), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_421), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_383), .B(n_360), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_384), .B(n_360), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g453 ( .A(n_406), .B(n_342), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_381), .B(n_357), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_384), .B(n_360), .Y(n_455) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_426), .A2(n_308), .A3(n_281), .B(n_366), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_385), .B(n_361), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_385), .B(n_361), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
OAI21xp33_ASAP7_75t_SL g460 ( .A1(n_406), .A2(n_353), .B(n_362), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_408), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_375), .B(n_337), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_374), .B(n_366), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_406), .A2(n_357), .B1(n_336), .B2(n_348), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_336), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_397), .B(n_336), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_411), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_374), .B(n_353), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_417), .B(n_353), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
NOR2x1p5_ASAP7_75t_L g474 ( .A(n_412), .B(n_348), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_417), .B(n_348), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_420), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_418), .B(n_348), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_382), .A2(n_362), .B(n_359), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_420), .Y(n_480) );
NOR2x1p5_ASAP7_75t_L g481 ( .A(n_412), .B(n_348), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_373), .Y(n_483) );
AND2x4_ASAP7_75t_SL g484 ( .A(n_387), .B(n_337), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_378), .B(n_337), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_418), .B(n_367), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
NAND2x1_ASAP7_75t_SL g489 ( .A(n_379), .B(n_367), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_379), .B(n_422), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_357), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_424), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_376), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_378), .B(n_341), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_422), .B(n_367), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_425), .Y(n_497) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_398), .A2(n_359), .B(n_357), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_376), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_425), .Y(n_500) );
AND2x4_ASAP7_75t_SL g501 ( .A(n_387), .B(n_341), .Y(n_501) );
AND3x2_ASAP7_75t_L g502 ( .A(n_405), .B(n_368), .C(n_341), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_372), .B(n_345), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_377), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_372), .B(n_345), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_431), .B(n_345), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_377), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_433), .B(n_351), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_434), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_428), .B(n_368), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_398), .B(n_351), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_400), .B(n_351), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_380), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_380), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_400), .B(n_368), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_405), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_456), .B(n_410), .C(n_386), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_483), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_436), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_490), .B(n_401), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_414), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_442), .B(n_447), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_460), .B(n_381), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_441), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_483), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_506), .B(n_427), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_516), .A2(n_399), .B(n_402), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_445), .B(n_432), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_503), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_443), .Y(n_531) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_489), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_448), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_505), .B(n_432), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_451), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_479), .A2(n_404), .B1(n_401), .B2(n_390), .C(n_392), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_474), .B(n_387), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_437), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_491), .B(n_414), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_439), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_471), .B(n_404), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_461), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_442), .B(n_388), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_467), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_471), .B(n_435), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_469), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_453), .B(n_466), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_511), .B(n_407), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_472), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_440), .B(n_465), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_473), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_481), .B(n_381), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_466), .B(n_381), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_463), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g562 ( .A1(n_498), .A2(n_409), .B(n_407), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_470), .B(n_409), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_447), .B(n_388), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_477), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_484), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_512), .B(n_434), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_480), .Y(n_568) );
OAI21xp33_ASAP7_75t_SL g569 ( .A1(n_450), .A2(n_389), .B(n_392), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_464), .A2(n_396), .B(n_394), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_470), .B(n_387), .Y(n_571) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_484), .B(n_391), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_450), .B(n_415), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_455), .B(n_389), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_457), .Y(n_575) );
NOR2xp67_ASAP7_75t_SL g576 ( .A(n_462), .B(n_391), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_482), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_487), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_455), .B(n_394), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_458), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_458), .B(n_396), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_488), .B(n_364), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_475), .B(n_364), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_475), .B(n_364), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_493), .B(n_364), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_496), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_478), .B(n_364), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_478), .B(n_314), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_572), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_517), .A2(n_515), .B1(n_454), .B2(n_486), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_553), .A2(n_502), .B(n_501), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_562), .A2(n_515), .B1(n_454), .B2(n_486), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_549), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
OAI311xp33_ASAP7_75t_L g599 ( .A1(n_537), .A2(n_494), .A3(n_485), .B1(n_508), .C1(n_514), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_571), .B(n_544), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_547), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_537), .B(n_510), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_569), .A2(n_513), .B1(n_507), .B2(n_504), .C(n_509), .Y(n_603) );
AO32x1_ASAP7_75t_L g604 ( .A1(n_566), .A2(n_501), .A3(n_444), .B1(n_497), .B2(n_500), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_564), .Y(n_606) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_558), .B(n_454), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_588), .B(n_510), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_523), .B(n_502), .C(n_500), .Y(n_609) );
OAI322xp33_ASAP7_75t_SL g610 ( .A1(n_520), .A2(n_495), .A3(n_446), .B1(n_444), .B2(n_438), .C1(n_497), .C2(n_17), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_588), .B(n_438), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_538), .A2(n_495), .B1(n_446), .B2(n_300), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_559), .A2(n_289), .B(n_311), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g615 ( .A1(n_573), .A2(n_314), .A3(n_291), .B1(n_287), .B2(n_15), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_520), .A2(n_311), .B(n_292), .Y(n_616) );
OAI322xp33_ASAP7_75t_L g617 ( .A1(n_574), .A2(n_11), .A3(n_12), .B1(n_13), .B2(n_16), .C1(n_18), .C2(n_19), .Y(n_617) );
AOI32xp33_ASAP7_75t_L g618 ( .A1(n_518), .A2(n_314), .A3(n_291), .B1(n_287), .B2(n_16), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_574), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_519), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_529), .B(n_304), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_527), .B(n_304), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_524), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_531), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_532), .A2(n_292), .B(n_291), .C(n_287), .Y(n_625) );
NAND2xp33_ASAP7_75t_L g626 ( .A(n_538), .B(n_19), .Y(n_626) );
AOI21xp33_ASAP7_75t_SL g627 ( .A1(n_525), .A2(n_20), .B(n_290), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_527), .B(n_304), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_532), .A2(n_290), .B(n_304), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_533), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_539), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_558), .A2(n_291), .B(n_20), .C(n_290), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_526), .B(n_288), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_570), .B(n_189), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_518), .A2(n_186), .B(n_23), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_534), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_536), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_525), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_626), .B(n_570), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_599), .A2(n_528), .B(n_522), .C(n_577), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_598), .Y(n_641) );
AOI322xp5_ASAP7_75t_L g642 ( .A1(n_602), .A2(n_521), .A3(n_556), .B1(n_563), .B2(n_542), .C1(n_575), .C2(n_581), .Y(n_642) );
NAND5xp2_ASAP7_75t_L g643 ( .A(n_595), .B(n_591), .C(n_586), .D(n_589), .E(n_585), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_594), .A2(n_530), .B1(n_576), .B2(n_580), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_607), .A2(n_550), .B(n_580), .C(n_540), .Y(n_645) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_603), .A2(n_590), .A3(n_557), .B(n_584), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_610), .A2(n_555), .B1(n_541), .B2(n_546), .C(n_579), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_601), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_596), .A2(n_582), .B1(n_560), .B2(n_543), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_606), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_593), .A2(n_551), .B1(n_548), .B2(n_578), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_604), .A2(n_577), .B(n_583), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_612), .B(n_561), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_619), .B(n_552), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_631), .B(n_554), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_593), .A2(n_535), .B1(n_567), .B2(n_568), .Y(n_656) );
OAI322xp33_ASAP7_75t_SL g657 ( .A1(n_592), .A2(n_587), .A3(n_583), .B1(n_565), .B2(n_288), .C1(n_32), .C2(n_33), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_604), .A2(n_587), .B(n_288), .Y(n_658) );
AOI321xp33_ASAP7_75t_L g659 ( .A1(n_613), .A2(n_288), .A3(n_27), .B1(n_29), .B2(n_30), .C(n_35), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_627), .A2(n_605), .B(n_617), .C(n_634), .Y(n_660) );
OAI322xp33_ASAP7_75t_L g661 ( .A1(n_638), .A2(n_186), .A3(n_288), .B1(n_36), .B2(n_39), .C1(n_40), .C2(n_41), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g662 ( .A1(n_609), .A2(n_22), .B(n_42), .C(n_45), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_632), .A2(n_280), .B(n_54), .C(n_56), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_597), .A2(n_280), .B1(n_62), .B2(n_63), .C(n_65), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_621), .A2(n_47), .B(n_66), .C(n_67), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_604), .A2(n_69), .B(n_70), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_616), .A2(n_71), .B(n_72), .C(n_74), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_622), .A2(n_75), .B1(n_76), .B2(n_77), .C1(n_78), .C2(n_79), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_628), .A2(n_82), .B1(n_83), .B2(n_85), .C1(n_86), .C2(n_87), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_620), .A2(n_89), .B1(n_92), .B2(n_94), .C(n_96), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_635), .B(n_98), .C(n_99), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_615), .B(n_100), .C(n_618), .D(n_608), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_623), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_624), .A2(n_630), .B1(n_636), .B2(n_637), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_625), .A2(n_614), .B(n_611), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_600), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_629), .A2(n_610), .B1(n_599), .B2(n_603), .C(n_602), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_655), .B(n_676), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_677), .B(n_639), .C(n_646), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_660), .B(n_642), .C(n_675), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_662), .B(n_643), .C(n_659), .D(n_668), .Y(n_681) );
AND4x1_ASAP7_75t_L g682 ( .A(n_669), .B(n_666), .C(n_640), .D(n_665), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_672), .A2(n_644), .B1(n_656), .B2(n_647), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_647), .B(n_674), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_684), .B(n_673), .Y(n_685) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_682), .B(n_671), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_678), .B(n_651), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_679), .Y(n_688) );
NOR3x2_ASAP7_75t_L g689 ( .A(n_686), .B(n_680), .C(n_683), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_688), .B(n_652), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_685), .B(n_681), .C(n_670), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_690), .B(n_687), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_689), .Y(n_693) );
OAI21x1_ASAP7_75t_L g694 ( .A1(n_692), .A2(n_685), .B(n_691), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_693), .A2(n_687), .B1(n_645), .B2(n_649), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_694), .A2(n_663), .B(n_650), .C(n_641), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_695), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_648), .B1(n_664), .B2(n_654), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_696), .B(n_657), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_667), .B(n_653), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_700), .A2(n_658), .B1(n_633), .B2(n_661), .Y(n_701) );
endmodule