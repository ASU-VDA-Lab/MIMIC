module real_jpeg_25934_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_33),
.B1(n_150),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_150),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_1),
.A2(n_71),
.B1(n_72),
.B2(n_150),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_10),
.B1(n_34),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_161),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_4),
.A2(n_71),
.B1(n_72),
.B2(n_161),
.Y(n_253)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_6),
.A2(n_115),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_24),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_158),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_67),
.C(n_72),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_52),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_6),
.A2(n_91),
.B1(n_247),
.B2(n_253),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_40),
.B1(n_71),
.B2(n_72),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_9),
.A2(n_58),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_9),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_140)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_34),
.B1(n_75),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_75),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_12),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_152),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_71),
.B1(n_72),
.B2(n_152),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_12),
.A2(n_114),
.B1(n_115),
.B2(n_152),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_14),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_35),
.B1(n_71),
.B2(n_72),
.Y(n_178)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_15),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_87),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_20),
.B(n_76),
.CI(n_87),
.CON(n_330),
.SN(n_330)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_21),
.A2(n_22),
.B1(n_110),
.B2(n_123),
.Y(n_109)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_47),
.C(n_62),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B(n_37),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_23),
.B(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_23),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_23),
.B(n_105),
.Y(n_307)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_24),
.A2(n_41),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_41),
.B1(n_160),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_24),
.A2(n_41),
.B1(n_168),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_25),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_25),
.A2(n_29),
.B(n_157),
.C(n_174),
.Y(n_173)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_25),
.B(n_158),
.CON(n_202),
.SN(n_202)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_26),
.B(n_28),
.C(n_106),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_26),
.A2(n_51),
.A3(n_54),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_29),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_31),
.Y(n_112)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_41),
.A2(n_104),
.B(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_41),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_41),
.A2(n_288),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_56),
.B(n_59),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_48),
.B(n_61),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_48),
.A2(n_52),
.B1(n_193),
.B2(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_50),
.B(n_53),
.Y(n_203)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_52),
.B(n_121),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_54),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_54),
.B(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_60),
.A2(n_78),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_62),
.A2(n_63),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B(n_73),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_74),
.B(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_65),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_65),
.A2(n_83),
.B(n_209),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_65),
.A2(n_208),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_65),
.A2(n_207),
.B1(n_208),
.B2(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_65),
.A2(n_100),
.B1(n_208),
.B2(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_86),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_84),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_70),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_70),
.B(n_158),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_71),
.B(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_76),
.A2(n_77),
.B(n_81),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_78),
.A2(n_80),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_78),
.A2(n_120),
.B(n_151),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_78),
.A2(n_80),
.B1(n_149),
.B2(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_79),
.A2(n_80),
.B(n_122),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_102),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_88),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_89),
.A2(n_90),
.B1(n_99),
.B2(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_89),
.A2(n_90),
.B1(n_102),
.B2(n_103),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B(n_97),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_91),
.A2(n_97),
.B(n_141),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_91),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_91),
.A2(n_244),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_92),
.A2(n_93),
.B1(n_140),
.B2(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_92),
.B(n_142),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_92),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_98),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_106),
.B(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_124),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_121),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_327),
.B(n_331),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_314),
.B(n_326),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_296),
.B(n_313),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_194),
.B(n_273),
.C(n_295),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_179),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_164),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_145),
.B1(n_162),
.B2(n_163),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_135),
.B(n_163),
.C(n_164),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_136),
.B(n_138),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_158),
.B(n_187),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_172),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_293)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_180),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_183),
.B(n_185),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_188),
.B(n_238),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_268),
.B(n_272),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_221),
.B(n_267),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_210),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_199),
.B(n_210),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_204),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_205),
.B(n_206),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_218),
.C(n_220),
.Y(n_269)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_262),
.B(n_266),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_240),
.B(n_261),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_249),
.B(n_260),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_248),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_255),
.B(n_259),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_275),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_293),
.B2(n_294),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_284),
.C(n_294),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_283),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_289),
.C(n_292),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_312),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_302),
.B1(n_310),
.B2(n_311),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_311),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_306),
.C(n_308),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_324),
.B2(n_325),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_323),
.C(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_329),
.B(n_330),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_330),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);


endmodule