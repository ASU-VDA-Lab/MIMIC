module fake_jpeg_21954_n_47 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_14),
.B1(n_13),
.B2(n_27),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_5),
.C(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_25),
.B2(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_14),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_29),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_R g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_9),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_11),
.Y(n_47)
);


endmodule