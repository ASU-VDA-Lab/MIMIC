module fake_jpeg_10346_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_33),
.B1(n_25),
.B2(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_64),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_48),
.B1(n_20),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_50),
.B1(n_51),
.B2(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_95),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_48),
.B1(n_31),
.B2(n_30),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_76),
.B1(n_25),
.B2(n_33),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_78),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_27),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_27),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_98),
.Y(n_120)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_92),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_63),
.B(n_32),
.Y(n_124)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_64),
.B(n_62),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_113),
.B(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_114),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_49),
.B1(n_57),
.B2(n_47),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_26),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_124),
.B1(n_32),
.B2(n_34),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_51),
.B1(n_47),
.B2(n_33),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_57),
.B1(n_25),
.B2(n_66),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_125),
.B1(n_26),
.B2(n_29),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_126),
.Y(n_142)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_133),
.Y(n_177)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_22),
.B(n_18),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_148),
.B1(n_156),
.B2(n_108),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_59),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_152),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_36),
.B1(n_117),
.B2(n_121),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_112),
.B1(n_109),
.B2(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_108),
.B1(n_101),
.B2(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_57),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_74),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_86),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_129),
.C(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_32),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_159),
.B(n_34),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_175),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_109),
.B1(n_110),
.B2(n_101),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_165),
.A2(n_180),
.B1(n_147),
.B2(n_154),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_109),
.B(n_118),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_176),
.B(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_SL g219 ( 
.A(n_167),
.B(n_170),
.C(n_174),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_172),
.C(n_182),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_129),
.B1(n_35),
.B2(n_78),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_186),
.B1(n_188),
.B2(n_157),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_148),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_118),
.B(n_40),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_38),
.B(n_34),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_22),
.B(n_18),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_141),
.B1(n_146),
.B2(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_193),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_40),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_130),
.A2(n_38),
.B(n_85),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_191),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_130),
.A2(n_35),
.B1(n_0),
.B2(n_2),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_35),
.B1(n_0),
.B2(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_0),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_1),
.C(n_3),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_197),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_201),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_142),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_132),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_213),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_150),
.B1(n_135),
.B2(n_151),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_215),
.B1(n_219),
.B2(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_133),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_220),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_133),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_164),
.B(n_175),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_SL g266 ( 
.A(n_225),
.B(n_235),
.C(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_168),
.C(n_171),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_238),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_170),
.B(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_239),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_180),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_188),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_174),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_191),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_175),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_169),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_169),
.B1(n_182),
.B2(n_179),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_223),
.B1(n_212),
.B2(n_195),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_267),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_225),
.B1(n_199),
.B2(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_262),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_205),
.B(n_214),
.C(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_234),
.B(n_232),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_245),
.B1(n_237),
.B2(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_222),
.C(n_224),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_271),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_209),
.B1(n_222),
.B2(n_169),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_1),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_202),
.B1(n_209),
.B2(n_194),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_240),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_242),
.Y(n_273)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_233),
.C(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_278),
.C(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_227),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_235),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_229),
.C(n_196),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_262),
.C(n_252),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_267),
.C(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_292),
.B(n_294),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_260),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_302),
.C(n_303),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_300),
.B1(n_276),
.B2(n_275),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_257),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_256),
.C(n_258),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_265),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_278),
.C(n_288),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_309),
.B(n_312),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_280),
.C(n_283),
.Y(n_309)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_4),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_299),
.B(n_296),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_5),
.C(n_6),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_7),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_7),
.C(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_314),
.B(n_316),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_297),
.B1(n_10),
.B2(n_11),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_306),
.B(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_9),
.Y(n_327)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_12),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_12),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_330),
.B(n_328),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_318),
.B(n_323),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.C(n_329),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.A3(n_324),
.B1(n_321),
.B2(n_317),
.C1(n_334),
.C2(n_15),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_13),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_13),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_14),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_14),
.B(n_326),
.Y(n_341)
);


endmodule