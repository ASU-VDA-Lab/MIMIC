module real_jpeg_4029_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx5_ASAP7_75t_L g186 ( 
.A(n_0),
.Y(n_186)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_0),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_1),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_1),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_2),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_2),
.A2(n_179),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_2),
.A2(n_108),
.B1(n_179),
.B2(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_2),
.A2(n_179),
.B1(n_324),
.B2(n_400),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_210),
.B1(n_229),
.B2(n_233),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_3),
.A2(n_100),
.B1(n_210),
.B2(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_3),
.A2(n_47),
.B1(n_210),
.B2(n_420),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_5),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_60),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_6),
.A2(n_60),
.B1(n_230),
.B2(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_6),
.A2(n_60),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_7),
.A2(n_95),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_7),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_162),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_7),
.A2(n_102),
.B1(n_162),
.B2(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_7),
.A2(n_162),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_12),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_12),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_124),
.C(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_12),
.B(n_90),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_12),
.B(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_166),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_12),
.B(n_103),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_13),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_14),
.A2(n_73),
.B1(n_221),
.B2(n_309),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_14),
.A2(n_73),
.B1(n_284),
.B2(n_387),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_14),
.A2(n_73),
.B1(n_396),
.B2(n_397),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_15),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_50),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_50),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_15),
.A2(n_50),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_17),
.A2(n_177),
.B1(n_229),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_17),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_17),
.A2(n_278),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_17),
.A2(n_278),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_278),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_18),
.A2(n_47),
.B1(n_54),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_18),
.A2(n_75),
.B1(n_130),
.B2(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_18),
.A2(n_75),
.B1(n_155),
.B2(n_366),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_18),
.A2(n_75),
.B1(n_266),
.B2(n_434),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_523),
.B(n_525),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_51),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_24),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_24),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_28),
.Y(n_323)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_29),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_29),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_32),
.Y(n_332)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_36),
.A2(n_348),
.B(n_351),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_36),
.B(n_353),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_39),
.Y(n_326)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_42),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_51)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_47),
.B(n_159),
.Y(n_333)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_51),
.B(n_65),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_61),
.B1(n_69),
.B2(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_52),
.A2(n_53),
.B1(n_61),
.B2(n_74),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_52),
.A2(n_352),
.B(n_399),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_52),
.A2(n_61),
.B1(n_399),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_52),
.A2(n_61),
.B1(n_69),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_58),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_61),
.B(n_159),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_61),
.A2(n_419),
.B(n_448),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_143),
.B(n_522),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_139),
.C(n_140),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_66),
.A2(n_67),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_76),
.C(n_112),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_68),
.B(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_76),
.A2(n_112),
.B1(n_113),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_76),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_77),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_77),
.A2(n_104),
.B1(n_299),
.B2(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_77),
.A2(n_104),
.B1(n_391),
.B2(n_395),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_77),
.A2(n_99),
.B1(n_104),
.B2(n_499),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_84),
.Y(n_363)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_87),
.Y(n_288)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_90),
.A2(n_141),
.B1(n_304),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_90),
.A2(n_141),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_90)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_93),
.Y(n_261)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_94),
.Y(n_407)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_96),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_96),
.Y(n_405)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_100),
.Y(n_435)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_104),
.B(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_104),
.A2(n_299),
.B(n_303),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_106),
.Y(n_394)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_108),
.Y(n_273)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_108),
.A2(n_260),
.A3(n_270),
.B1(n_280),
.B2(n_283),
.Y(n_279)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_111),
.Y(n_268)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_111),
.Y(n_393)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_111),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_112),
.A2(n_113),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_112),
.B(n_494),
.C(n_497),
.Y(n_505)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_126),
.B(n_135),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_153),
.B(n_160),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_114),
.A2(n_126),
.B1(n_207),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_114),
.A2(n_160),
.B(n_259),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_114),
.A2(n_126),
.B1(n_365),
.B2(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_115),
.B(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_115),
.A2(n_166),
.B1(n_386),
.B2(n_388),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_115),
.A2(n_166),
.B1(n_388),
.B2(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_115),
.A2(n_166),
.B1(n_404),
.B2(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_119),
.Y(n_262)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_207),
.B(n_214),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_126),
.A2(n_214),
.B(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_134),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_134),
.Y(n_383)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_135),
.Y(n_438)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_138),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_139),
.B(n_140),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_141),
.A2(n_265),
.B(n_271),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_141),
.B(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_141),
.A2(n_271),
.B(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_516),
.B(n_521),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_488),
.B(n_513),
.Y(n_144)
);

OAI311xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_372),
.A3(n_464),
.B1(n_482),
.C1(n_487),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_314),
.B(n_371),
.Y(n_146)
);

AO21x1_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_290),
.B(n_313),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_253),
.B(n_289),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_217),
.B(n_252),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_173),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_151),
.B(n_173),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_167),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_152),
.A2(n_167),
.B1(n_168),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_156),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_156),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_159),
.A2(n_184),
.B(n_191),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g265 ( 
.A1(n_159),
.A2(n_266),
.B(n_269),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_159),
.A2(n_333),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_204),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_205),
.C(n_216),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_184),
.B(n_191),
.Y(n_174)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_184),
.A2(n_336),
.B1(n_337),
.B2(n_339),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_184),
.A2(n_247),
.B1(n_378),
.B2(n_382),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_184),
.A2(n_193),
.B(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_195),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_185),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_185),
.A2(n_277),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_185),
.A2(n_340),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_197),
.Y(n_309)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_215),
.B2(n_216),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_241),
.B(n_251),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_240),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_239),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_239),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_238),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_247),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_249),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_247),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_255),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_274),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_263),
.B2(n_264),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_263),
.C(n_274),
.Y(n_291)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_291),
.B(n_292),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_312),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_296),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_306),
.C(n_307),
.Y(n_342)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_315),
.B(n_316),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_345),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_317)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_334),
.B2(n_335),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_320),
.B(n_334),
.Y(n_459)
);

OAI32xp33_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_324),
.A3(n_326),
.B1(n_327),
.B2(n_333),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_342),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_342),
.B(n_343),
.C(n_345),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_358),
.B2(n_370),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_346),
.B(n_359),
.C(n_364),
.Y(n_473)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_358),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_364),
.Y(n_358)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_449),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_373),
.A2(n_449),
.B(n_483),
.C(n_486),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_425),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_374),
.B(n_425),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_401),
.C(n_410),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_401),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_389),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_390),
.C(n_398),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_385),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_385),
.Y(n_455)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_398),
.Y(n_389)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

INVx8_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_408),
.B2(n_409),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_408),
.Y(n_442)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_408),
.A2(n_409),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_408),
.A2(n_442),
.B(n_445),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.C(n_423),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_414),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_417),
.A2(n_418),
.B1(n_423),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_426),
.B(n_429),
.C(n_440),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_440),
.B2(n_441),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_436),
.B(n_439),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_437),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_439),
.B(n_491),
.CI(n_492),
.CON(n_490),
.SN(n_490)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_491),
.C(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_462),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_462),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_455),
.C(n_456),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_452),
.B1(n_455),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_455),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_475),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.C(n_460),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_477),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_474),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_474),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_471),
.C(n_473),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_480),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_471),
.A2(n_472),
.B1(n_473),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_479),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_502),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_501),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_501),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_490),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_496),
.B2(n_500),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_494),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_504),
.C(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_512),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_512),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_520),
.Y(n_521)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx13_ASAP7_75t_L g527 ( 
.A(n_524),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_528),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);


endmodule