module fake_jpeg_5578_n_189 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_37),
.B1(n_22),
.B2(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_46),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_22),
.B1(n_15),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_70),
.B1(n_76),
.B2(n_35),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_55),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_64),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_47),
.B(n_42),
.C(n_45),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_53),
.B(n_70),
.C(n_76),
.Y(n_87)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_33),
.A2(n_37),
.B1(n_26),
.B2(n_20),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_15),
.B(n_30),
.C(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_72),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_20),
.B1(n_31),
.B2(n_21),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_73),
.C(n_11),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_31),
.B1(n_21),
.B2(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_32),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_29),
.C(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_4),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_24),
.B1(n_14),
.B2(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_34),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_35),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_88),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_100),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_59),
.B1(n_65),
.B2(n_62),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_7),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_8),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_12),
.B(n_11),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_97),
.C(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_56),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_90),
.B1(n_81),
.B2(n_101),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_123),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_60),
.B1(n_75),
.B2(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_49),
.B1(n_48),
.B2(n_69),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_48),
.B(n_64),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_73),
.B1(n_51),
.B2(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_52),
.B1(n_79),
.B2(n_12),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_86),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_11),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_91),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_93),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_113),
.B(n_86),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_80),
.B1(n_96),
.B2(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_105),
.B1(n_123),
.B2(n_111),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_135),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_122),
.C(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_90),
.B1(n_81),
.B2(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_120),
.B(n_122),
.Y(n_145)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_112),
.C(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_141),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_128),
.A3(n_136),
.B1(n_137),
.B2(n_149),
.C1(n_130),
.C2(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_153),
.C(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_131),
.B(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_131),
.B1(n_130),
.B2(n_132),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_105),
.B1(n_117),
.B2(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_125),
.B(n_52),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_159),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_164),
.B(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_166),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_116),
.C(n_129),
.Y(n_166)
);

AO221x1_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_138),
.B1(n_133),
.B2(n_134),
.C(n_100),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_157),
.B1(n_161),
.B2(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_148),
.B1(n_156),
.B2(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_146),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_95),
.C(n_85),
.Y(n_179)
);

AOI222xp33_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_165),
.B1(n_145),
.B2(n_166),
.C1(n_141),
.C2(n_84),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_177),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_89),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_91),
.B1(n_85),
.B2(n_79),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_174),
.C(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_176),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_182),
.B(n_95),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);


endmodule