module fake_aes_5537_n_524 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_524);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_524;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g74 ( .A(n_1), .Y(n_74) );
BUFx6f_ASAP7_75t_L g75 ( .A(n_27), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_6), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_34), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_11), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_33), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_36), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_66), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_11), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_4), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_53), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_29), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_0), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_30), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_58), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_1), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_56), .Y(n_101) );
BUFx10_ASAP7_75t_L g102 ( .A(n_44), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_73), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_16), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_51), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_26), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_95), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_102), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_96), .B(n_0), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_84), .B(n_2), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
AND2x6_ASAP7_75t_L g121 ( .A(n_95), .B(n_28), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_74), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_75), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_102), .B(n_3), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_101), .B(n_5), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_97), .B(n_5), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_112), .B(n_102), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_117), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_112), .B(n_103), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_112), .B(n_102), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_112), .B(n_76), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_117), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_115), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_115), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_117), .B(n_76), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
INVx5_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_124), .B(n_77), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_130), .Y(n_151) );
BUFx10_ASAP7_75t_L g152 ( .A(n_121), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_124), .B(n_81), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_130), .B(n_87), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_128), .B(n_82), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_155), .A2(n_130), .B1(n_121), .B2(n_131), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_149), .B(n_118), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_139), .B(n_128), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_136), .B(n_118), .Y(n_164) );
OR2x6_ASAP7_75t_L g165 ( .A(n_151), .B(n_122), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_151), .B(n_126), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_155), .A2(n_121), .B1(n_133), .B2(n_131), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_139), .B(n_122), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_136), .B(n_133), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_155), .A2(n_129), .B1(n_98), .B2(n_78), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_147), .A2(n_144), .B(n_157), .C(n_159), .Y(n_178) );
INVxp67_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_147), .B(n_92), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
AND3x1_ASAP7_75t_SL g183 ( .A(n_155), .B(n_86), .C(n_105), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_138), .B(n_86), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_155), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_121), .B1(n_88), .B2(n_105), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_178), .A2(n_134), .B(n_150), .C(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_168), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_174), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_174), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_164), .B(n_155), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_192), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_177), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_177), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_188), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_185), .B(n_149), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_192), .B(n_149), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_156), .B(n_100), .C(n_88), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_180), .A2(n_149), .B(n_132), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_185), .B(n_149), .Y(n_209) );
AOI22xp33_ASAP7_75t_SL g210 ( .A1(n_165), .A2(n_108), .B1(n_146), .B2(n_121), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_182), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_146), .B1(n_121), .B2(n_111), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_184), .B(n_152), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_188), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_161), .A2(n_123), .B1(n_100), .B2(n_111), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_188), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
CKINVDCx8_ASAP7_75t_R g220 ( .A(n_186), .Y(n_220) );
BUFx2_ASAP7_75t_SL g221 ( .A(n_175), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_184), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g225 ( .A1(n_219), .A2(n_172), .B1(n_176), .B2(n_166), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_219), .A2(n_172), .B1(n_184), .B2(n_166), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_219), .B(n_166), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_223), .B(n_163), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_208), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_208), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_222), .A2(n_181), .B1(n_191), .B2(n_179), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_222), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_210), .A2(n_171), .B1(n_181), .B2(n_170), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_199), .B(n_223), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_196), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_199), .B(n_175), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_196), .B(n_175), .Y(n_238) );
INVx4_ASAP7_75t_L g239 ( .A(n_211), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_220), .B(n_175), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_222), .A2(n_189), .B1(n_167), .B2(n_170), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_189), .B1(n_162), .B2(n_190), .Y(n_244) );
OAI221xp5_ASAP7_75t_L g245 ( .A1(n_198), .A2(n_183), .B1(n_123), .B2(n_89), .C(n_104), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_220), .B(n_175), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_190), .B1(n_132), .B2(n_93), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_221), .B(n_187), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_197), .A2(n_132), .B1(n_169), .B2(n_175), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_240), .B(n_197), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_240), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_233), .B(n_201), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_217), .B1(n_195), .B2(n_200), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_249), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_201), .B(n_204), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_239), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_225), .A2(n_217), .B1(n_200), .B2(n_215), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_215), .B1(n_213), .B2(n_204), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_233), .B(n_201), .Y(n_261) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_206), .B(n_193), .C(n_204), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g263 ( .A1(n_230), .A2(n_212), .B1(n_221), .B2(n_214), .Y(n_263) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_228), .A2(n_212), .B1(n_209), .B2(n_218), .C(n_216), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_246), .Y(n_265) );
OAI21xp33_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_234), .B(n_248), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_212), .B1(n_218), .B2(n_216), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_209), .B1(n_202), .B2(n_224), .C(n_91), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_202), .B1(n_203), .B2(n_224), .Y(n_270) );
OAI31xp33_ASAP7_75t_L g271 ( .A1(n_242), .A2(n_87), .A3(n_91), .B(n_93), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_239), .B(n_203), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_250), .B(n_224), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_250), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_268), .Y(n_275) );
AOI33xp33_ASAP7_75t_L g276 ( .A1(n_255), .A2(n_94), .A3(n_99), .B1(n_104), .B2(n_106), .B3(n_107), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_265), .B(n_227), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_269), .A2(n_235), .B1(n_227), .B2(n_232), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_269), .A2(n_227), .B1(n_232), .B2(n_235), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_266), .A2(n_235), .B1(n_202), .B2(n_243), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_254), .B(n_202), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_268), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_266), .A2(n_238), .B1(n_237), .B2(n_249), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
OAI21xp33_ASAP7_75t_SL g286 ( .A1(n_254), .A2(n_239), .B(n_249), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_271), .B(n_79), .C(n_99), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_238), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_261), .B(n_238), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_274), .B(n_238), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_265), .Y(n_292) );
OAI211xp5_ASAP7_75t_SL g293 ( .A1(n_271), .A2(n_94), .B(n_106), .C(n_107), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_274), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_256), .B(n_249), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_259), .A2(n_244), .B1(n_109), .B2(n_207), .C(n_241), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_274), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_279), .A2(n_264), .B1(n_262), .B2(n_260), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_283), .B(n_252), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_277), .B(n_256), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_286), .A2(n_264), .B(n_263), .C(n_272), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_289), .B(n_261), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_286), .A2(n_257), .B(n_265), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_283), .B(n_252), .Y(n_306) );
OAI33xp33_ASAP7_75t_L g307 ( .A1(n_279), .A2(n_109), .A3(n_110), .B1(n_114), .B2(n_113), .B3(n_127), .Y(n_307) );
AOI31xp33_ASAP7_75t_L g308 ( .A1(n_280), .A2(n_263), .A3(n_267), .B(n_270), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_275), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_290), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_252), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_290), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_294), .B(n_253), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_262), .A3(n_261), .B(n_253), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_110), .B1(n_257), .B2(n_273), .C(n_79), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
OAI31xp33_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_273), .A3(n_251), .B(n_203), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_295), .A2(n_272), .B1(n_258), .B2(n_237), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_276), .B(n_127), .C(n_119), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_292), .B(n_278), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_284), .B(n_127), .C(n_119), .D(n_114), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_291), .B(n_258), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_311), .B(n_278), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_318), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_304), .B(n_277), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_301), .B(n_295), .Y(n_334) );
NOR3xp33_ASAP7_75t_SL g335 ( .A(n_302), .B(n_296), .C(n_83), .Y(n_335) );
NOR2xp67_ASAP7_75t_L g336 ( .A(n_305), .B(n_277), .Y(n_336) );
NOR2x1_ASAP7_75t_L g337 ( .A(n_309), .B(n_288), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_327), .B(n_288), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_320), .B(n_277), .Y(n_340) );
OAI22xp33_ASAP7_75t_SL g341 ( .A1(n_299), .A2(n_288), .B1(n_295), .B2(n_282), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_308), .A2(n_295), .B1(n_281), .B2(n_258), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_324), .B(n_258), .Y(n_343) );
OAI21xp33_ASAP7_75t_SL g344 ( .A1(n_299), .A2(n_247), .B(n_258), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_307), .A2(n_258), .B1(n_79), .B2(n_237), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_322), .B(n_79), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_7), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_326), .B(n_7), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_312), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_312), .B(n_79), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_300), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_301), .B(n_326), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_306), .B(n_79), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_301), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_306), .B(n_113), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_303), .B(n_113), .Y(n_362) );
AND3x2_ASAP7_75t_L g363 ( .A(n_319), .B(n_8), .C(n_9), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_298), .B(n_114), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_301), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_321), .B(n_119), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_125), .B1(n_140), .B2(n_207), .C(n_158), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_316), .B(n_125), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_325), .B(n_9), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_317), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_304), .B(n_125), .Y(n_371) );
NAND2xp33_ASAP7_75t_SL g372 ( .A(n_331), .B(n_237), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_328), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_345), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_330), .B(n_10), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_349), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_357), .B(n_10), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_352), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_356), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_343), .Y(n_383) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_337), .B(n_125), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_125), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_355), .B(n_12), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_336), .A2(n_140), .B(n_203), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_365), .B(n_13), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_332), .B(n_13), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_360), .B(n_14), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_332), .B(n_14), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_351), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_348), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_343), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_340), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_360), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_341), .A2(n_140), .B1(n_158), .B2(n_148), .C(n_141), .Y(n_400) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_371), .B(n_211), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_358), .B(n_333), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_338), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_344), .B(n_15), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_329), .B(n_15), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_358), .B(n_16), .Y(n_406) );
AOI31xp33_ASAP7_75t_L g407 ( .A1(n_342), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_354), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_350), .B(n_17), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_350), .B(n_211), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_361), .B(n_18), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_334), .B(n_20), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_364), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_334), .B(n_21), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_372), .A2(n_369), .B(n_346), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_403), .B(n_370), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_394), .B(n_364), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_399), .B(n_368), .Y(n_420) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_391), .B(n_335), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_398), .B(n_363), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_373), .B(n_368), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_407), .A2(n_369), .B1(n_366), .B2(n_367), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_393), .B(n_22), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_383), .B(n_23), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_397), .B(n_24), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_380), .A2(n_158), .B(n_148), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_372), .A2(n_211), .B1(n_158), .B2(n_148), .Y(n_432) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_404), .B(n_211), .Y(n_433) );
XOR2x2_ASAP7_75t_L g434 ( .A(n_406), .B(n_25), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
AOI322xp5_ASAP7_75t_L g436 ( .A1(n_377), .A2(n_31), .A3(n_32), .B1(n_35), .B2(n_37), .C1(n_38), .C2(n_39), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_408), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_377), .B(n_187), .C(n_41), .D(n_46), .Y(n_438) );
XOR2xp5_ASAP7_75t_L g439 ( .A(n_405), .B(n_40), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_416), .B(n_47), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_379), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_390), .B(n_48), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_390), .B(n_49), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_387), .A2(n_205), .B1(n_54), .B2(n_55), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_402), .B(n_52), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_385), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_381), .B(n_60), .Y(n_452) );
AOI21xp33_ASAP7_75t_SL g453 ( .A1(n_391), .A2(n_61), .B(n_62), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_392), .B(n_382), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_391), .B(n_148), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
AOI32xp33_ASAP7_75t_L g457 ( .A1(n_386), .A2(n_63), .A3(n_69), .B1(n_71), .B2(n_187), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_392), .B(n_141), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_411), .A2(n_141), .B1(n_143), .B2(n_145), .C(n_148), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_401), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_414), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_395), .B(n_141), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_386), .A2(n_141), .B(n_143), .C(n_145), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
AOI322xp5_ASAP7_75t_L g466 ( .A1(n_389), .A2(n_141), .A3(n_143), .B1(n_145), .B2(n_148), .C1(n_158), .C2(n_205), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_400), .A2(n_143), .B(n_145), .C(n_158), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_396), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_415), .A2(n_205), .B1(n_145), .B2(n_143), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_412), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_389), .B(n_143), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_412), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_415), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_388), .A2(n_169), .B1(n_342), .B2(n_372), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_388), .A2(n_169), .B1(n_342), .B2(n_372), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_403), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_403), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_403), .B(n_394), .Y(n_479) );
XOR2x2_ASAP7_75t_L g480 ( .A(n_406), .B(n_379), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_404), .B(n_399), .Y(n_481) );
BUFx8_ASAP7_75t_L g482 ( .A(n_446), .Y(n_482) );
OAI211xp5_ASAP7_75t_L g483 ( .A1(n_421), .A2(n_481), .B(n_422), .C(n_447), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_418), .B(n_442), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_438), .B(n_433), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_447), .A2(n_437), .B1(n_472), .B2(n_470), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_480), .A2(n_442), .B(n_479), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g488 ( .A1(n_457), .A2(n_459), .B(n_440), .C(n_458), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_440), .A2(n_476), .B1(n_474), .B2(n_455), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_435), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_455), .A2(n_434), .B(n_417), .Y(n_492) );
OAI22x1_ASAP7_75t_L g493 ( .A1(n_439), .A2(n_473), .B1(n_448), .B2(n_460), .Y(n_493) );
NAND3xp33_ASAP7_75t_SL g494 ( .A(n_453), .B(n_463), .C(n_431), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_464), .B(n_469), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_478), .B(n_477), .Y(n_496) );
AOI31xp33_ASAP7_75t_L g497 ( .A1(n_425), .A2(n_445), .A3(n_448), .B(n_443), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_424), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_445), .A2(n_454), .B(n_469), .C(n_444), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_467), .B(n_436), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_483), .B(n_420), .C(n_467), .D(n_423), .Y(n_501) );
XOR2x2_ASAP7_75t_L g502 ( .A(n_486), .B(n_419), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_487), .A2(n_461), .B1(n_468), .B2(n_465), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_497), .A2(n_450), .B1(n_449), .B2(n_464), .Y(n_504) );
AO22x2_ASAP7_75t_L g505 ( .A1(n_489), .A2(n_428), .B1(n_429), .B2(n_475), .Y(n_505) );
OAI211xp5_ASAP7_75t_L g506 ( .A1(n_499), .A2(n_466), .B(n_432), .C(n_427), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_491), .Y(n_507) );
INVxp33_ASAP7_75t_L g508 ( .A(n_493), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_490), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_508), .A2(n_484), .B1(n_485), .B2(n_495), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_507), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_503), .A2(n_496), .B1(n_498), .B2(n_450), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_509), .Y(n_513) );
NAND3xp33_ASAP7_75t_SL g514 ( .A(n_500), .B(n_488), .C(n_430), .Y(n_514) );
OAI222xp33_ASAP7_75t_L g515 ( .A1(n_510), .A2(n_504), .B1(n_501), .B2(n_505), .C1(n_502), .C2(n_506), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_511), .A2(n_505), .B1(n_451), .B2(n_456), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_513), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_516), .A2(n_514), .B1(n_512), .B2(n_494), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_517), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_518), .A2(n_515), .B1(n_482), .B2(n_452), .Y(n_520) );
XNOR2xp5_ASAP7_75t_L g521 ( .A(n_519), .B(n_482), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_521), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_522), .A2(n_520), .B(n_426), .C(n_441), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_523), .A2(n_471), .B(n_462), .Y(n_524) );
endmodule