module real_aes_17086_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g109 ( .A(n_0), .B(n_110), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_1), .A2(n_34), .B1(n_154), .B2(n_246), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_2), .A2(n_9), .B1(n_551), .B2(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_4), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_5), .A2(n_10), .B1(n_552), .B2(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g117 ( .A(n_6), .B(n_30), .Y(n_117) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_7), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_8), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_11), .B(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_12), .A2(n_99), .B1(n_199), .B2(n_551), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_13), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_14), .A2(n_31), .B1(n_569), .B2(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_15), .B(n_169), .Y(n_566) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_16), .A2(n_48), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_17), .B(n_250), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_18), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_19), .A2(n_39), .B1(n_206), .B2(n_221), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_20), .Y(n_274) );
INVx1_ASAP7_75t_L g873 ( .A(n_21), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_22), .A2(n_45), .B1(n_221), .B2(n_551), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_23), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_24), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_25), .B(n_229), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_26), .Y(n_558) );
XNOR2x1_ASAP7_75t_L g129 ( .A(n_27), .B(n_40), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_28), .B(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_29), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_32), .A2(n_84), .B1(n_154), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_33), .A2(n_37), .B1(n_154), .B2(n_554), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_35), .A2(n_51), .B1(n_551), .B2(n_606), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_36), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_38), .Y(n_865) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_41), .B(n_169), .Y(n_217) );
INVx2_ASAP7_75t_L g123 ( .A(n_42), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_43), .B(n_202), .Y(n_244) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
BUFx3_ASAP7_75t_L g126 ( .A(n_44), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_46), .B(n_188), .Y(n_252) );
XOR2x2_ASAP7_75t_L g136 ( .A(n_47), .B(n_137), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_47), .A2(n_858), .B1(n_859), .B2(n_862), .Y(n_857) );
INVx1_ASAP7_75t_L g862 ( .A(n_47), .Y(n_862) );
AND2x2_ASAP7_75t_L g280 ( .A(n_49), .B(n_188), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_50), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_52), .B(n_229), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_53), .B(n_206), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_54), .A2(n_71), .B1(n_206), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_55), .A2(n_74), .B1(n_154), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_56), .B(n_310), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_57), .A2(n_158), .B(n_167), .C(n_273), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_58), .A2(n_96), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
AND2x4_ASAP7_75t_L g172 ( .A(n_60), .B(n_173), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_61), .A2(n_62), .B1(n_221), .B2(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_63), .A2(n_81), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_63), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_64), .B(n_147), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_65), .B(n_188), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_66), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_67), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g173 ( .A(n_68), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_69), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_70), .B(n_147), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_72), .B(n_154), .Y(n_305) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_73), .B(n_202), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_75), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g160 ( .A(n_76), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_77), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_78), .B(n_169), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_79), .B(n_163), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_80), .A2(n_95), .B1(n_167), .B2(n_221), .Y(n_538) );
INVx1_ASAP7_75t_L g861 ( .A(n_81), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_82), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_83), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_85), .A2(n_90), .B1(n_228), .B2(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_86), .B(n_169), .Y(n_201) );
NAND2xp33_ASAP7_75t_SL g186 ( .A(n_87), .B(n_157), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_88), .B(n_200), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_89), .B(n_147), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_91), .Y(n_591) );
INVx1_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_92), .B(n_844), .Y(n_843) );
NAND2xp33_ASAP7_75t_L g570 ( .A(n_93), .B(n_169), .Y(n_570) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_94), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_97), .B(n_188), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_98), .B(n_157), .C(n_181), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_100), .B(n_154), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_101), .B(n_229), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_118), .B(n_872), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx12f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_SL g876 ( .A(n_106), .Y(n_876) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_115), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .C(n_113), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AND3x2_ASAP7_75t_L g854 ( .A(n_111), .B(n_113), .C(n_127), .Y(n_854) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g844 ( .A(n_112), .Y(n_844) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g127 ( .A(n_117), .Y(n_127) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_117), .B(n_126), .Y(n_871) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_836), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_128), .Y(n_119) );
BUFx12f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_L g850 ( .A(n_123), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_123), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_SL g842 ( .A(n_127), .B(n_843), .Y(n_842) );
XOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AOI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .B(n_525), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g525 ( .A(n_132), .B(n_526), .Y(n_525) );
INVx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx12f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g870 ( .A(n_135), .B(n_871), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_137), .A2(n_856), .B1(n_857), .B2(n_863), .Y(n_855) );
INVx2_ASAP7_75t_L g863 ( .A(n_137), .Y(n_863) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_457), .Y(n_137) );
NAND4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_332), .C(n_372), .D(n_421), .Y(n_138) );
NOR2xp67_ASAP7_75t_L g139 ( .A(n_140), .B(n_281), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_191), .B1(n_253), .B2(n_262), .Y(n_140) );
INVx1_ASAP7_75t_L g453 ( .A(n_141), .Y(n_453) );
INVx1_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_142), .B(n_300), .Y(n_369) );
AND2x2_ASAP7_75t_L g400 ( .A(n_142), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_174), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_143), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g324 ( .A(n_143), .Y(n_324) );
AND2x2_ASAP7_75t_L g499 ( .A(n_143), .B(n_367), .Y(n_499) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx2_ASAP7_75t_L g264 ( .A(n_144), .Y(n_264) );
AND2x2_ASAP7_75t_L g352 ( .A(n_144), .B(n_314), .Y(n_352) );
AND2x2_ASAP7_75t_L g396 ( .A(n_144), .B(n_301), .Y(n_396) );
OR2x2_ASAP7_75t_L g414 ( .A(n_144), .B(n_415), .Y(n_414) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g318 ( .A(n_145), .B(n_301), .Y(n_318) );
BUFx2_ASAP7_75t_L g375 ( .A(n_145), .Y(n_375) );
OR2x2_ASAP7_75t_L g383 ( .A(n_145), .B(n_341), .Y(n_383) );
INVx1_ASAP7_75t_L g438 ( .A(n_145), .Y(n_438) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_L g578 ( .A(n_147), .Y(n_578) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_SL g170 ( .A(n_148), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_SL g177 ( .A(n_148), .Y(n_177) );
INVx2_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
BUFx3_ASAP7_75t_L g534 ( .A(n_148), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_148), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g562 ( .A(n_148), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_148), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_148), .B(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_161), .B(n_170), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_158), .Y(n_152) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_154), .A2(n_221), .B1(n_278), .B2(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g552 ( .A(n_154), .Y(n_552) );
INVx4_ASAP7_75t_L g554 ( .A(n_154), .Y(n_554) );
INVx1_ASAP7_75t_L g606 ( .A(n_154), .Y(n_606) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_155), .Y(n_157) );
INVx1_ASAP7_75t_L g167 ( .A(n_155), .Y(n_167) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_155), .Y(n_169) );
INVx1_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
INVx1_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_155), .Y(n_221) );
INVx1_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_155), .Y(n_246) );
INVx2_ASAP7_75t_L g275 ( .A(n_155), .Y(n_275) );
INVx2_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
INVx1_ASAP7_75t_L g569 ( .A(n_157), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_158), .A2(n_184), .B(n_186), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_158), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_158), .A2(n_305), .B(n_306), .Y(n_304) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g165 ( .A(n_160), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
BUFx8_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B1(n_166), .B2(n_168), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_163), .A2(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_169), .A2(n_180), .B(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
INVx3_ASAP7_75t_L g551 ( .A(n_169), .Y(n_551) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_171), .A2(n_179), .B(n_183), .Y(n_178) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_171), .A2(n_197), .B(n_203), .Y(n_196) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_171), .A2(n_215), .B(n_218), .Y(n_214) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_171), .A2(n_243), .B(n_247), .Y(n_242) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_171), .A2(n_304), .B(n_307), .Y(n_303) );
BUFx10_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx10_ASAP7_75t_L g237 ( .A(n_172), .Y(n_237) );
INVx1_ASAP7_75t_L g541 ( .A(n_172), .Y(n_541) );
AND2x2_ASAP7_75t_L g265 ( .A(n_174), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g377 ( .A(n_174), .B(n_354), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_174), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g415 ( .A(n_175), .Y(n_415) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_175), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_175), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g327 ( .A(n_176), .B(n_267), .Y(n_327) );
INVx1_ASAP7_75t_L g341 ( .A(n_176), .Y(n_341) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_187), .Y(n_176) );
INVx1_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
INVx1_ASAP7_75t_L g539 ( .A(n_181), .Y(n_539) );
INVx1_ASAP7_75t_SL g555 ( .A(n_181), .Y(n_555) );
INVx1_ASAP7_75t_L g597 ( .A(n_185), .Y(n_597) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g195 ( .A(n_189), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_189), .B(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_189), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g236 ( .A(n_190), .Y(n_236) );
INVx2_ASAP7_75t_L g240 ( .A(n_190), .Y(n_240) );
NAND2x1_ASAP7_75t_L g191 ( .A(n_192), .B(n_208), .Y(n_191) );
AND2x4_ASAP7_75t_L g502 ( .A(n_192), .B(n_430), .Y(n_502) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_193), .Y(n_261) );
BUFx3_ASAP7_75t_L g296 ( .A(n_193), .Y(n_296) );
INVx1_ASAP7_75t_L g362 ( .A(n_193), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_193), .B(n_211), .Y(n_365) );
AND2x2_ASAP7_75t_L g390 ( .A(n_193), .B(n_241), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_193), .Y(n_393) );
AND2x2_ASAP7_75t_L g425 ( .A(n_193), .B(n_290), .Y(n_425) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_207), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_195), .A2(n_196), .B(n_207), .Y(n_291) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_195), .A2(n_303), .B(n_312), .Y(n_302) );
OAI21xp33_ASAP7_75t_SL g330 ( .A1(n_195), .A2(n_303), .B(n_312), .Y(n_330) );
O2A1O1Ixp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_201), .C(n_202), .Y(n_197) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_202), .A2(n_219), .B(n_220), .Y(n_218) );
INVx6_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g564 ( .A1(n_202), .A2(n_554), .B(n_565), .C(n_566), .Y(n_564) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_223), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g334 ( .A(n_210), .B(n_320), .Y(n_334) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g360 ( .A(n_212), .B(n_347), .Y(n_360) );
AND2x2_ASAP7_75t_L g389 ( .A(n_212), .B(n_225), .Y(n_389) );
OR2x2_ASAP7_75t_L g485 ( .A(n_212), .B(n_225), .Y(n_485) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_222), .Y(n_212) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_242), .B(n_252), .Y(n_241) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_213), .A2(n_214), .B(n_222), .Y(n_259) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_213), .A2(n_242), .B(n_252), .Y(n_290) );
INVx2_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_221), .A2(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g364 ( .A(n_223), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g513 ( .A(n_223), .Y(n_513) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
OR2x2_ASAP7_75t_L g447 ( .A(n_224), .B(n_257), .Y(n_447) );
INVx1_ASAP7_75t_L g469 ( .A(n_224), .Y(n_469) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_241), .Y(n_224) );
AND2x2_ASAP7_75t_L g285 ( .A(n_225), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g320 ( .A(n_225), .B(n_290), .Y(n_320) );
INVx1_ASAP7_75t_L g347 ( .A(n_225), .Y(n_347) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_225), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_225), .B(n_241), .Y(n_434) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_236), .A3(n_237), .B(n_238), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_231), .B1(n_232), .B2(n_234), .Y(n_226) );
INVx1_ASAP7_75t_L g588 ( .A(n_229), .Y(n_588) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_231), .A2(n_536), .B1(n_538), .B2(n_539), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_231), .A2(n_550), .B1(n_553), .B2(n_555), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_231), .A2(n_568), .B(n_570), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_231), .A2(n_234), .B1(n_576), .B2(n_577), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_231), .A2(n_555), .B1(n_587), .B2(n_589), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_231), .A2(n_234), .B1(n_596), .B2(n_598), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_231), .A2(n_234), .B1(n_605), .B2(n_607), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_231), .A2(n_234), .B1(n_621), .B2(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g599 ( .A(n_233), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_234), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
INVx2_ASAP7_75t_L g269 ( .A(n_236), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_236), .B(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_236), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g270 ( .A(n_237), .Y(n_270) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_237), .A2(n_575), .A3(n_578), .B(n_579), .Y(n_574) );
AO31x2_ASAP7_75t_L g585 ( .A1(n_237), .A2(n_548), .A3(n_586), .B(n_590), .Y(n_585) );
AO31x2_ASAP7_75t_L g594 ( .A1(n_237), .A2(n_534), .A3(n_595), .B(n_600), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
BUFx2_ASAP7_75t_L g548 ( .A(n_240), .Y(n_548) );
AND2x2_ASAP7_75t_L g371 ( .A(n_241), .B(n_291), .Y(n_371) );
INVx2_ASAP7_75t_L g310 ( .A(n_246), .Y(n_310) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_251), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR3x1_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .C(n_260), .Y(n_254) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_257), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g319 ( .A(n_257), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g370 ( .A(n_257), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g410 ( .A(n_257), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_257), .B(n_433), .Y(n_465) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_258), .B(n_346), .Y(n_406) );
AND2x2_ASAP7_75t_L g430 ( .A(n_258), .B(n_290), .Y(n_430) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g286 ( .A(n_259), .Y(n_286) );
BUFx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g441 ( .A(n_261), .B(n_320), .Y(n_441) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_264), .B(n_327), .Y(n_506) );
AND2x4_ASAP7_75t_L g498 ( .A(n_265), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_265), .B(n_318), .Y(n_512) );
INVx2_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
INVx2_ASAP7_75t_L g402 ( .A(n_266), .Y(n_402) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g386 ( .A(n_267), .Y(n_386) );
AOI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_280), .Y(n_267) );
NOR2xp67_ASAP7_75t_SL g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g603 ( .A(n_269), .Y(n_603) );
INVx1_ASAP7_75t_L g556 ( .A(n_270), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_SL g537 ( .A(n_275), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_321), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_297), .B1(n_315), .B2(n_319), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_292), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g349 ( .A(n_285), .B(n_296), .Y(n_349) );
AND2x2_ASAP7_75t_L g509 ( .A(n_285), .B(n_390), .Y(n_509) );
BUFx2_ASAP7_75t_L g380 ( .A(n_286), .Y(n_380) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g379 ( .A(n_289), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g294 ( .A(n_290), .Y(n_294) );
INVx1_ASAP7_75t_L g346 ( .A(n_290), .Y(n_346) );
INVx1_ASAP7_75t_L g471 ( .A(n_291), .Y(n_471) );
AOI31xp33_ASAP7_75t_L g489 ( .A1(n_292), .A2(n_490), .A3(n_491), .B(n_492), .Y(n_489) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_294), .B(n_389), .Y(n_488) );
INVx2_ASAP7_75t_L g516 ( .A(n_294), .Y(n_516) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_295), .Y(n_331) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g344 ( .A(n_296), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_296), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g474 ( .A(n_296), .B(n_434), .Y(n_474) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_313), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g385 ( .A(n_301), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_311), .Y(n_307) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
INVx1_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
AND2x2_ASAP7_75t_L g419 ( .A(n_318), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g475 ( .A(n_318), .B(n_402), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_319), .A2(n_392), .B(n_394), .Y(n_391) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_331), .Y(n_321) );
NAND3x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .C(n_328), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g493 ( .A(n_324), .B(n_413), .Y(n_493) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NOR2x1_ASAP7_75t_SL g446 ( .A(n_326), .B(n_358), .Y(n_446) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g366 ( .A(n_327), .B(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_328), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_328), .B(n_437), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_328), .B(n_437), .Y(n_510) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g413 ( .A(n_330), .B(n_386), .Y(n_413) );
AND2x2_ASAP7_75t_L g333 ( .A(n_331), .B(n_334), .Y(n_333) );
AOI221x1_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B1(n_342), .B2(n_351), .C(n_355), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g514 ( .A1(n_334), .A2(n_515), .A3(n_520), .B1(n_521), .B2(n_523), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_339), .B(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
OR2x2_ASAP7_75t_L g470 ( .A(n_341), .B(n_471), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_348), .C(n_350), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g392 ( .A(n_345), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g409 ( .A(n_345), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_348), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_444) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g522 ( .A(n_352), .Y(n_522) );
INVx2_ASAP7_75t_L g367 ( .A(n_354), .Y(n_367) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_363), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g491 ( .A(n_360), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_361), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B1(n_368), .B2(n_370), .Y(n_363) );
AND2x4_ASAP7_75t_L g460 ( .A(n_366), .B(n_375), .Y(n_460) );
INVx1_ASAP7_75t_L g519 ( .A(n_367), .Y(n_519) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g398 ( .A(n_371), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_371), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_371), .B(n_399), .Y(n_490) );
AOI211x1_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_379), .B(n_381), .C(n_407), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR3x2_ASAP7_75t_L g482 ( .A(n_375), .B(n_377), .C(n_378), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_398), .B1(n_400), .B2(n_403), .Y(n_397) );
NOR2x1p5_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_377), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
INVx2_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_387), .B(n_391), .C(n_397), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_389), .B(n_393), .Y(n_404) );
INVx1_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_389), .B(n_496), .Y(n_504) );
OAI32xp33_ASAP7_75t_L g479 ( .A1(n_390), .A2(n_435), .A3(n_480), .B1(n_482), .B2(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g496 ( .A(n_390), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_390), .B(n_410), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_393), .B(n_427), .Y(n_462) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g440 ( .A(n_399), .B(n_425), .Y(n_440) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g449 ( .A(n_402), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g417 ( .A(n_405), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B1(n_416), .B2(n_418), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g436 ( .A(n_413), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_413), .B(n_420), .Y(n_524) );
INVx1_ASAP7_75t_SL g450 ( .A(n_414), .Y(n_450) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_444), .C(n_451), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_435), .B(n_439), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_428), .Y(n_423) );
INVxp67_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g481 ( .A(n_426), .Y(n_481) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .C(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g443 ( .A(n_437), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g452 ( .A(n_440), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_445), .A2(n_496), .B1(n_497), .B2(n_500), .C(n_501), .Y(n_495) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI32xp33_ASAP7_75t_L g451 ( .A1(n_448), .A2(n_452), .A3(n_453), .B1(n_454), .B2(n_456), .Y(n_451) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_454), .A2(n_464), .B1(n_465), .B2(n_466), .C(n_472), .Y(n_463) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_476), .C(n_494), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B(n_463), .Y(n_458) );
AOI211x1_ASAP7_75t_L g476 ( .A1(n_459), .A2(n_477), .B(n_479), .C(n_486), .Y(n_476) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2x1_ASAP7_75t_SL g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g478 ( .A(n_469), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AO21x1_ASAP7_75t_L g486 ( .A1(n_475), .A2(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g520 ( .A(n_491), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI21xp33_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_511), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g517 ( .A(n_516), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND4xp75_ASAP7_75t_L g526 ( .A(n_527), .B(n_676), .C(n_752), .D(n_804), .Y(n_526) );
AND3x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_649), .C(n_662), .Y(n_527) );
AOI221x1_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_581), .B1(n_610), .B2(n_614), .C(n_626), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_529), .A2(n_650), .B(n_652), .C(n_653), .Y(n_649) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_544), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g613 ( .A(n_533), .Y(n_613) );
BUFx2_ASAP7_75t_L g631 ( .A(n_533), .Y(n_631) );
OR2x2_ASAP7_75t_L g673 ( .A(n_533), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g680 ( .A(n_533), .B(n_547), .Y(n_680) );
AND2x4_ASAP7_75t_L g715 ( .A(n_533), .B(n_546), .Y(n_715) );
OR2x2_ASAP7_75t_L g758 ( .A(n_533), .B(n_574), .Y(n_758) );
AO31x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .A3(n_540), .B(n_542), .Y(n_533) );
AO31x2_ASAP7_75t_L g602 ( .A1(n_540), .A2(n_603), .A3(n_604), .B(n_608), .Y(n_602) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g571 ( .A(n_541), .Y(n_571) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_559), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_546), .B(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_546), .Y(n_645) );
INVx2_ASAP7_75t_L g672 ( .A(n_546), .Y(n_672) );
INVx3_ASAP7_75t_L g685 ( .A(n_546), .Y(n_685) );
AND2x2_ASAP7_75t_L g803 ( .A(n_546), .B(n_632), .Y(n_803) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g612 ( .A(n_547), .B(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .A3(n_556), .B(n_557), .Y(n_547) );
AO31x2_ASAP7_75t_L g619 ( .A1(n_556), .A2(n_603), .A3(n_620), .B(n_623), .Y(n_619) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g688 ( .A(n_560), .Y(n_688) );
INVx1_ASAP7_75t_L g815 ( .A(n_560), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_573), .Y(n_560) );
AND2x2_ASAP7_75t_L g611 ( .A(n_561), .B(n_574), .Y(n_611) );
INVx1_ASAP7_75t_L g674 ( .A(n_561), .Y(n_674) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_572), .Y(n_561) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_562), .A2(n_563), .B(n_572), .Y(n_633) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_567), .B(n_571), .Y(n_563) );
INVx2_ASAP7_75t_L g629 ( .A(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g681 ( .A(n_573), .B(n_632), .Y(n_681) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_574), .Y(n_703) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_583), .A2(n_675), .B1(n_679), .B2(n_682), .Y(n_678) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_592), .Y(n_583) );
INVx1_ASAP7_75t_L g696 ( .A(n_584), .Y(n_696) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g616 ( .A(n_585), .B(n_594), .Y(n_616) );
AND2x2_ASAP7_75t_L g647 ( .A(n_585), .B(n_602), .Y(n_647) );
INVx4_ASAP7_75t_SL g658 ( .A(n_585), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_585), .B(n_692), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_585), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_707), .Y(n_729) );
OR2x2_ASAP7_75t_L g762 ( .A(n_593), .B(n_744), .Y(n_762) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_602), .Y(n_593) );
INVx2_ASAP7_75t_L g636 ( .A(n_594), .Y(n_636) );
INVx1_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
AND2x2_ASAP7_75t_L g648 ( .A(n_594), .B(n_618), .Y(n_648) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_594), .Y(n_664) );
INVx1_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_594), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g625 ( .A(n_602), .Y(n_625) );
AND2x4_ASAP7_75t_L g635 ( .A(n_602), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g661 ( .A(n_602), .Y(n_661) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_602), .Y(n_738) );
INVx1_ASAP7_75t_L g831 ( .A(n_602), .Y(n_831) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_611), .B(n_684), .Y(n_751) );
AND2x2_ASAP7_75t_L g764 ( .A(n_611), .B(n_680), .Y(n_764) );
AND2x2_ASAP7_75t_L g834 ( .A(n_611), .B(n_685), .Y(n_834) );
AND2x4_ASAP7_75t_L g669 ( .A(n_613), .B(n_632), .Y(n_669) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g736 ( .A(n_616), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g750 ( .A(n_616), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_616), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g652 ( .A(n_617), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_617), .B(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g746 ( .A1(n_617), .A2(n_747), .B(n_750), .C(n_751), .Y(n_746) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_625), .Y(n_617) );
AND2x2_ASAP7_75t_L g717 ( .A(n_618), .B(n_658), .Y(n_717) );
INVx3_ASAP7_75t_L g744 ( .A(n_618), .Y(n_744) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g639 ( .A(n_619), .Y(n_639) );
AND2x4_ASAP7_75t_L g665 ( .A(n_619), .B(n_625), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_625), .B(n_658), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_634), .B1(n_642), .B2(n_646), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g783 ( .A(n_628), .Y(n_783) );
AND2x4_ASAP7_75t_L g694 ( .A(n_629), .B(n_674), .Y(n_694) );
INVx1_ASAP7_75t_L g714 ( .A(n_629), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_631), .A2(n_687), .B1(n_697), .B2(n_699), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_631), .B(n_688), .Y(n_745) );
NAND2x1_ASAP7_75t_L g802 ( .A(n_631), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g817 ( .A(n_631), .Y(n_817) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g756 ( .A(n_633), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
AND2x2_ASAP7_75t_L g675 ( .A(n_635), .B(n_657), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_635), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g716 ( .A(n_635), .B(n_717), .Y(n_716) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_635), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_635), .B(n_698), .Y(n_797) );
AND2x4_ASAP7_75t_L g820 ( .A(n_635), .B(n_748), .Y(n_820) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx3_ASAP7_75t_L g698 ( .A(n_638), .Y(n_698) );
AND2x2_ASAP7_75t_L g710 ( .A(n_638), .B(n_703), .Y(n_710) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g660 ( .A(n_639), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g708 ( .A(n_639), .Y(n_708) );
INVx1_ASAP7_75t_L g651 ( .A(n_640), .Y(n_651) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g808 ( .A(n_641), .B(n_658), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g734 ( .A(n_643), .B(n_715), .Y(n_734) );
INVx2_ASAP7_75t_L g775 ( .A(n_643), .Y(n_775) );
AND2x4_ASAP7_75t_L g776 ( .A(n_643), .B(n_669), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_644), .B(n_694), .Y(n_824) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_647), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g719 ( .A(n_647), .B(n_664), .Y(n_719) );
INVx1_ASAP7_75t_L g811 ( .A(n_647), .Y(n_811) );
AND2x2_ASAP7_75t_L g810 ( .A(n_648), .B(n_737), .Y(n_810) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_652), .A2(n_782), .B1(n_784), .B2(n_786), .Y(n_781) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g690 ( .A(n_658), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g726 ( .A(n_658), .Y(n_726) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_658), .Y(n_732) );
INVx2_ASAP7_75t_L g749 ( .A(n_658), .Y(n_749) );
OR2x2_ASAP7_75t_L g770 ( .A(n_658), .B(n_733), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_658), .B(n_728), .Y(n_780) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g747 ( .A(n_660), .B(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_660), .Y(n_801) );
INVx1_ASAP7_75t_L g728 ( .A(n_661), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_670), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_665), .B(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g733 ( .A(n_665), .Y(n_733) );
AND2x2_ASAP7_75t_L g807 ( .A(n_665), .B(n_808), .Y(n_807) );
AOI211x1_ASAP7_75t_SL g735 ( .A1(n_666), .A2(n_736), .B(n_739), .C(n_746), .Y(n_735) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g792 ( .A(n_668), .B(n_669), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_669), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_669), .Y(n_785) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g700 ( .A(n_672), .Y(n_700) );
NOR2x1p5_ASAP7_75t_L g757 ( .A(n_672), .B(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_673), .B(n_702), .Y(n_701) );
NOR2xp67_ASAP7_75t_SL g774 ( .A(n_673), .B(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_L g835 ( .A(n_675), .B(n_743), .Y(n_835) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_720), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_686), .C(n_704), .Y(n_677) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_680), .Y(n_711) );
AND2x2_ASAP7_75t_L g718 ( .A(n_680), .B(n_714), .Y(n_718) );
AND2x4_ASAP7_75t_SL g832 ( .A(n_680), .B(n_694), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_681), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_683), .A2(n_725), .B1(n_797), .B2(n_798), .Y(n_796) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_L g814 ( .A(n_685), .B(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_693), .B2(n_695), .Y(n_687) );
NAND2x1_ASAP7_75t_L g763 ( .A(n_690), .B(n_743), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_690), .B(n_737), .Y(n_773) );
INVx1_ASAP7_75t_L g800 ( .A(n_690), .Y(n_800) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_693), .A2(n_819), .B(n_822), .Y(n_818) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_694), .A2(n_706), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g779 ( .A(n_698), .Y(n_779) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g723 ( .A(n_701), .Y(n_723) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_711), .B1(n_712), .B2(n_716), .C1(n_718), .C2(n_719), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g739 ( .A1(n_706), .A2(n_740), .B(n_745), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_707), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g821 ( .A(n_707), .Y(n_821) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_708), .Y(n_827) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
AND2x2_ASAP7_75t_L g791 ( .A(n_713), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g784 ( .A(n_714), .B(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_735), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_730), .B2(n_734), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_729), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g741 ( .A(n_727), .Y(n_741) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g769 ( .A(n_744), .B(n_761), .Y(n_769) );
OR2x2_ASAP7_75t_L g829 ( .A(n_744), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND5xp2_ASAP7_75t_L g805 ( .A(n_750), .B(n_797), .C(n_806), .D(n_809), .E(n_811), .Y(n_805) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_788), .Y(n_752) );
NAND2xp67_ASAP7_75t_SL g753 ( .A(n_754), .B(n_771), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_759), .B1(n_764), .B2(n_765), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NAND3xp33_ASAP7_75t_SL g759 ( .A(n_760), .B(n_762), .C(n_763), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g794 ( .A(n_763), .Y(n_794) );
NAND3xp33_ASAP7_75t_SL g765 ( .A(n_766), .B(n_769), .C(n_770), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g787 ( .A(n_768), .Y(n_787) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_769), .A2(n_800), .B(n_801), .C(n_802), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B1(n_776), .B2(n_777), .C(n_781), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_778), .B(n_826), .Y(n_825) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g795 ( .A(n_782), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_793), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g798 ( .A(n_792), .Y(n_798) );
AOI211xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_795), .B(n_796), .C(n_799), .Y(n_793) );
AOI211x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_812), .B(n_818), .C(n_833), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2x1p5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2x1_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_825), .B1(n_828), .B2(n_832), .Y(n_822) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_846), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_837), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_SL g838 ( .A(n_839), .B(n_845), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
CKINVDCx8_ASAP7_75t_R g841 ( .A(n_842), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_851), .B(n_864), .Y(n_846) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
CKINVDCx11_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
INVx4_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx10_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx4_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx4_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
endmodule