module fake_jpeg_24750_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_8),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_58),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_25),
.B1(n_18),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_63),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_46),
.B1(n_29),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_77),
.B1(n_90),
.B2(n_29),
.Y(n_108)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_71),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_29),
.B1(n_43),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_85),
.B1(n_97),
.B2(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_74),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_32),
.B1(n_63),
.B2(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_23),
.B(n_29),
.C(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_32),
.B1(n_43),
.B2(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_37),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_37),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_25),
.B1(n_35),
.B2(n_17),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_103),
.B1(n_111),
.B2(n_129),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_76),
.B1(n_95),
.B2(n_82),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_32),
.B1(n_45),
.B2(n_42),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_110),
.B1(n_119),
.B2(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_35),
.B1(n_17),
.B2(n_24),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_48),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_48),
.C(n_40),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_39),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_36),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_21),
.B(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_97),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_1),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_125),
.B(n_17),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_8),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_14),
.C(n_16),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_1),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_48),
.B1(n_40),
.B2(n_39),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_40),
.B1(n_39),
.B2(n_30),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_151),
.B1(n_28),
.B2(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_39),
.B1(n_40),
.B2(n_88),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_141),
.B1(n_124),
.B2(n_113),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_145),
.B(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_104),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_142),
.B1(n_156),
.B2(n_106),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_149),
.B(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_85),
.B1(n_95),
.B2(n_82),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_30),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_33),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_154),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_1),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_30),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_132),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_35),
.B(n_24),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_31),
.B(n_28),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

AO21x2_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_21),
.B(n_27),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_109),
.B(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_171),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_101),
.B1(n_115),
.B2(n_108),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_168),
.B1(n_155),
.B2(n_135),
.Y(n_192)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_150),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_118),
.B1(n_128),
.B2(n_110),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_128),
.C(n_119),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_135),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_120),
.B(n_123),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_184),
.B(n_125),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_112),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_145),
.Y(n_197)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_139),
.B(n_125),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_155),
.B(n_153),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_187),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_200),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_193),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_170),
.B1(n_178),
.B2(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_208),
.C(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_209),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_146),
.B(n_131),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_151),
.B1(n_145),
.B2(n_122),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_33),
.B1(n_34),
.B2(n_19),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_105),
.B(n_107),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_157),
.B(n_33),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_126),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_214),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_180),
.A2(n_126),
.B(n_129),
.C(n_116),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_217),
.B(n_28),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_159),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_171),
.A2(n_129),
.B(n_116),
.C(n_19),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_218),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_129),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_21),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_186),
.B1(n_176),
.B2(n_168),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_227),
.B1(n_233),
.B2(n_235),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_184),
.C(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_184),
.C(n_170),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_236),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_188),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_158),
.B1(n_113),
.B2(n_106),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_225),
.B1(n_202),
.B2(n_210),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_162),
.B1(n_116),
.B2(n_19),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_191),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_200),
.B1(n_189),
.B2(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_116),
.B(n_34),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_21),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_202),
.B1(n_194),
.B2(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_236),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_265),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_196),
.B(n_197),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_263),
.B(n_217),
.Y(n_279)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_196),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_223),
.B1(n_245),
.B2(n_239),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_243),
.B1(n_230),
.B2(n_234),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_229),
.B(n_215),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_222),
.B1(n_242),
.B2(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_224),
.C(n_226),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_277),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_244),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_243),
.B1(n_217),
.B2(n_212),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_254),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_235),
.B1(n_212),
.B2(n_219),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_252),
.B(n_247),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_217),
.B1(n_212),
.B2(n_27),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_212),
.CI(n_21),
.CON(n_284),
.SN(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_252),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_296),
.B1(n_284),
.B2(n_2),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_259),
.B1(n_272),
.B2(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_27),
.B1(n_3),
.B2(n_1),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_248),
.B(n_255),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_268),
.B(n_276),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_271),
.C(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_251),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_27),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_292),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_273),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_296),
.C(n_285),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_288),
.B1(n_297),
.B2(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_284),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_9),
.B(n_4),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_300),
.C(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_3),
.C(n_4),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_308),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_318),
.A2(n_320),
.B1(n_9),
.B2(n_4),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_287),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_301),
.B1(n_307),
.B2(n_5),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.C(n_11),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_313),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_11),
.Y(n_327)
);

OAI21x1_ASAP7_75t_SL g329 ( 
.A1(n_327),
.A2(n_11),
.B(n_5),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_325),
.B(n_315),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.C(n_330),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_327),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_324),
.B(n_331),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_323),
.A3(n_322),
.B1(n_7),
.B2(n_8),
.C1(n_13),
.C2(n_15),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_6),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_13),
.Y(n_337)
);

AOI311xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_13),
.A3(n_15),
.B(n_16),
.C(n_3),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_3),
.Y(n_339)
);


endmodule