module fake_jpeg_27596_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_31),
.B1(n_32),
.B2(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_41),
.B1(n_29),
.B2(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_54),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_19),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_30),
.C(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_27),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_71),
.Y(n_92)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_78),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_35),
.B1(n_41),
.B2(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_82),
.B1(n_85),
.B2(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_83),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_59),
.B1(n_57),
.B2(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_40),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_46),
.B1(n_52),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_93),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_54),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_57),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_38),
.C(n_72),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_54),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_38),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_67),
.B1(n_76),
.B2(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_126),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_95),
.B1(n_106),
.B2(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_116),
.Y(n_135)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_119),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_63),
.B(n_73),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_129),
.B(n_99),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_76),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_84),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_22),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_66),
.B(n_1),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_85),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_87),
.C(n_69),
.D(n_79),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_25),
.B(n_22),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_104),
.B1(n_81),
.B2(n_88),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_141),
.B(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_142),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_146),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_92),
.B(n_102),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_103),
.A3(n_15),
.B1(n_14),
.B2(n_12),
.C1(n_11),
.C2(n_9),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_92),
.B(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_111),
.A3(n_129),
.B1(n_118),
.B2(n_127),
.C1(n_119),
.C2(n_121),
.Y(n_155)
);

HAxp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_0),
.CON(n_146),
.SN(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_148),
.B(n_122),
.C(n_123),
.D(n_109),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_15),
.A3(n_14),
.B1(n_12),
.B2(n_9),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_117),
.C(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_159),
.C(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_161),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_162),
.C(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_114),
.C(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_169),
.C(n_149),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_153),
.B1(n_152),
.B2(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_151),
.C(n_159),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_137),
.CI(n_141),
.CON(n_174),
.SN(n_174)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_140),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_176),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_147),
.C(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_151),
.C(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_181),
.B(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_167),
.B1(n_166),
.B2(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_172),
.B1(n_170),
.B2(n_174),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_176),
.A3(n_146),
.B1(n_109),
.B2(n_120),
.C1(n_4),
.C2(n_0),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_1),
.C(n_3),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_160),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_120),
.B(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_185),
.B1(n_188),
.B2(n_6),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_195),
.B(n_4),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_185),
.B(n_8),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_3),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_191),
.B1(n_186),
.B2(n_8),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

AOI31xp33_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_199),
.A3(n_200),
.B(n_6),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_6),
.Y(n_203)
);


endmodule