module fake_ariane_2350_n_1639 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1639);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1639;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_60),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_80),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_96),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_99),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_19),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_35),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_44),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_74),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_69),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_45),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_26),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_17),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_29),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_37),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_90),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_20),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_78),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_11),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_46),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_147),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_15),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_0),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_46),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_101),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_64),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_51),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_106),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_84),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_26),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_89),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_92),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_63),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_71),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_154),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_102),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_43),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_150),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_105),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_95),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_130),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_125),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_86),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_44),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_10),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_13),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_30),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_14),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_1),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_139),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_123),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_65),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_116),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_134),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_54),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_34),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_23),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_9),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_67),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_53),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_12),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_122),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_94),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_81),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_132),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_11),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_141),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_42),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_72),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_163),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_76),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_160),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_100),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_129),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_62),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_104),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_53),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_126),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_6),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_38),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_128),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_49),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_83),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_108),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_42),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_66),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_219),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_R g328 ( 
.A(n_254),
.B(n_151),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_255),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_207),
.B(n_1),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_224),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_219),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_219),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_219),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_172),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_236),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_244),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_263),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_189),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_286),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_216),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_235),
.B(n_2),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_179),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_255),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_270),
.B(n_7),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_257),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_176),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_176),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_206),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_164),
.B(n_9),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_273),
.B(n_12),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_273),
.B(n_14),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_258),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_211),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_236),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_16),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_181),
.B(n_18),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_212),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_195),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_234),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_221),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_223),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_234),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_301),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_226),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_301),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_182),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_205),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_182),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_227),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_215),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_228),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_229),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_166),
.B(n_18),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_238),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_237),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_190),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_233),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_167),
.B(n_20),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_265),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_241),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_284),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_292),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_248),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_245),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_260),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_262),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_276),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_290),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_299),
.B(n_21),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_258),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_335),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_329),
.B(n_258),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_347),
.B(n_200),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_338),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_339),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_356),
.B(n_201),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_341),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_343),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_345),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_348),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_334),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_363),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_170),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_370),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_371),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_373),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_374),
.B(n_203),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_377),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_369),
.B(n_210),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_210),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_342),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_383),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_386),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_329),
.B(n_212),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_372),
.B(n_311),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_387),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_391),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_396),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_399),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_362),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_185),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_378),
.B(n_311),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_389),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_385),
.B(n_213),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_395),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_365),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_367),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_350),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_351),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_408),
.Y(n_483)
);

AO22x2_ASAP7_75t_L g484 ( 
.A1(n_407),
.A2(n_358),
.B1(n_397),
.B2(n_352),
.Y(n_484)
);

INVxp67_ASAP7_75t_R g485 ( 
.A(n_419),
.Y(n_485)
);

NAND2x1p5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_392),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_415),
.B(n_357),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_L g488 ( 
.A1(n_444),
.A2(n_353),
.B1(n_362),
.B2(n_354),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_340),
.Y(n_489)
);

BUFx8_ASAP7_75t_SL g490 ( 
.A(n_474),
.Y(n_490)
);

BUFx10_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_411),
.B(n_353),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_415),
.B(n_184),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_379),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_366),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_421),
.B(n_193),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_440),
.B(n_388),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_479),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_421),
.B(n_196),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_417),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_474),
.Y(n_513)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_466),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_459),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_464),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_394),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_433),
.B(n_340),
.C(n_330),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_407),
.B(n_393),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_437),
.B(n_202),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_407),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_328),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_441),
.B(n_346),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_471),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_448),
.B(n_393),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_448),
.B(n_406),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_441),
.B(n_448),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_465),
.B(n_318),
.Y(n_543)
);

AOI21x1_ASAP7_75t_L g544 ( 
.A1(n_430),
.A2(n_209),
.B(n_208),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_473),
.B(n_400),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_473),
.B(n_400),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_437),
.B(n_214),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_446),
.B(n_218),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_412),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_455),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_430),
.B(n_401),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_451),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_449),
.B(n_401),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_449),
.B(n_406),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_382),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_413),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_420),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_452),
.B(n_225),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_403),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_457),
.B(n_192),
.C(n_305),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_465),
.B(n_246),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_467),
.B(n_403),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_478),
.B(n_404),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_416),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_404),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_416),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_478),
.B(n_402),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_461),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_418),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_433),
.B(n_360),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_368),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_462),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_458),
.B(n_460),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_468),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_468),
.B(n_368),
.Y(n_582)
);

AO22x2_ASAP7_75t_L g583 ( 
.A1(n_468),
.A2(n_316),
.B1(n_320),
.B2(n_324),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_409),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_469),
.B(n_197),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_469),
.B(n_165),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_470),
.B(n_405),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_470),
.B(n_405),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_470),
.B(n_360),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_418),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_425),
.A2(n_361),
.B1(n_443),
.B2(n_454),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_422),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_425),
.B(n_239),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_432),
.B(n_251),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_409),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_409),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_423),
.B(n_261),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_432),
.B(n_165),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_434),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_414),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_414),
.B(n_361),
.Y(n_602)
);

NAND2x1p5_ASAP7_75t_L g603 ( 
.A(n_434),
.B(n_256),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_438),
.A2(n_312),
.B(n_295),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_426),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_438),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_414),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_443),
.B(n_169),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_168),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_442),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_447),
.B(n_281),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_454),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_442),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_SL g614 ( 
.A(n_463),
.B(n_185),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_466),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_472),
.B(n_398),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_450),
.B(n_169),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_584),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_486),
.B(n_171),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_486),
.B(n_171),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_522),
.A2(n_252),
.B1(n_323),
.B2(n_322),
.Y(n_623)
);

NOR2x1_ASAP7_75t_L g624 ( 
.A(n_498),
.B(n_289),
.Y(n_624)
);

OAI21xp33_ASAP7_75t_L g625 ( 
.A1(n_598),
.A2(n_303),
.B(n_192),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_522),
.B(n_173),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_571),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_499),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_489),
.B(n_431),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_519),
.A2(n_243),
.B(n_303),
.C(n_191),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_506),
.B(n_173),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_517),
.A2(n_243),
.B1(n_305),
.B2(n_186),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_504),
.B(n_174),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_489),
.B(n_186),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_481),
.A2(n_315),
.B(n_453),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_317),
.C(n_191),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_519),
.A2(n_604),
.B(n_501),
.C(n_540),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_542),
.A2(n_252),
.B1(n_323),
.B2(n_322),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_584),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_540),
.B(n_174),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_531),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_542),
.B(n_317),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_541),
.B(n_554),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_596),
.Y(n_644)
);

O2A1O1Ixp5_ASAP7_75t_L g645 ( 
.A1(n_539),
.A2(n_453),
.B(n_450),
.C(n_319),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_541),
.B(n_175),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_532),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_565),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_497),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_499),
.A2(n_321),
.B1(n_264),
.B2(n_253),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_175),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_583),
.A2(n_256),
.B1(n_259),
.B2(n_287),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_494),
.B(n_272),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_498),
.B(n_259),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_596),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_550),
.B(n_274),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_492),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_542),
.B(n_577),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_558),
.B(n_177),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_542),
.B(n_321),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_558),
.B(n_177),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_542),
.B(n_577),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_178),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_535),
.B(n_287),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_487),
.A2(n_198),
.B1(n_319),
.B2(n_313),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_499),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_583),
.A2(n_453),
.B1(n_450),
.B2(n_297),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_538),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_550),
.B(n_282),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_582),
.B(n_180),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_283),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_551),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_180),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_601),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_553),
.Y(n_677)
);

NOR3x1_ASAP7_75t_L g678 ( 
.A(n_566),
.B(n_293),
.C(n_294),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_601),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_589),
.B(n_183),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_561),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_183),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_574),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_487),
.A2(n_313),
.B1(n_308),
.B2(n_307),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_580),
.A2(n_296),
.B1(n_307),
.B2(n_306),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_573),
.B(n_536),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_570),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_573),
.B(n_187),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_308),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_588),
.B(n_306),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_574),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_588),
.B(n_304),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_513),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_575),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_574),
.Y(n_697)
);

BUFx6f_ASAP7_75t_SL g698 ( 
.A(n_535),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_499),
.A2(n_188),
.B1(n_300),
.B2(n_194),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_593),
.B(n_188),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_515),
.B(n_199),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_485),
.B(n_199),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_482),
.B(n_198),
.C(n_300),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_605),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_581),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_558),
.B(n_194),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_616),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_591),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_482),
.A2(n_249),
.B1(n_298),
.B2(n_288),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_563),
.B(n_25),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_513),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_602),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_543),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_516),
.B(n_217),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_581),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_495),
.B(n_29),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_529),
.B(n_32),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_32),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_607),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_520),
.B(n_222),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_557),
.B(n_33),
.Y(n_722)
);

CKINVDCx11_ASAP7_75t_R g723 ( 
.A(n_491),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_607),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_600),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_523),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_607),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_525),
.B(n_285),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_610),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_488),
.A2(n_250),
.B1(n_271),
.B2(n_269),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_610),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_526),
.B(n_230),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_528),
.B(n_231),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_530),
.B(n_232),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_543),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_491),
.B(n_36),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_557),
.B(n_247),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_612),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_492),
.Y(n_740)
);

BUFx8_ASAP7_75t_L g741 ( 
.A(n_490),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_557),
.B(n_266),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_610),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_503),
.A2(n_267),
.B(n_268),
.C(n_302),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_545),
.B(n_37),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_560),
.B(n_302),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_483),
.B(n_512),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_546),
.B(n_39),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_491),
.B(n_39),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_567),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_585),
.B(n_268),
.Y(n_751)
);

OAI21xp33_ASAP7_75t_L g752 ( 
.A1(n_599),
.A2(n_268),
.B(n_242),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_524),
.B(n_40),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_500),
.B(n_505),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_524),
.B(n_555),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_500),
.A2(n_268),
.B1(n_242),
.B2(n_168),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_41),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_555),
.B(n_41),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_555),
.B(n_47),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_493),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_560),
.B(n_268),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_585),
.B(n_47),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_505),
.B(n_48),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_585),
.B(n_48),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_490),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_496),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_592),
.B(n_49),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_641),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_629),
.B(n_512),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_637),
.A2(n_632),
.B(n_700),
.C(n_643),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_650),
.B(n_562),
.Y(n_771)
);

AOI21xp33_ASAP7_75t_L g772 ( 
.A1(n_763),
.A2(n_583),
.B(n_521),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_637),
.A2(n_502),
.B(n_511),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_647),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_658),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_700),
.A2(n_587),
.B(n_510),
.C(n_548),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_659),
.A2(n_509),
.B(n_507),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_711),
.A2(n_552),
.B(n_533),
.C(n_547),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_634),
.B(n_615),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_704),
.B(n_576),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_618),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_662),
.A2(n_511),
.B(n_502),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_657),
.A2(n_484),
.B1(n_614),
.B2(n_602),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_549),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_687),
.A2(n_484),
.B1(n_547),
.B2(n_508),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_669),
.Y(n_786)
);

AO21x1_ASAP7_75t_L g787 ( 
.A1(n_763),
.A2(n_613),
.B(n_539),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_736),
.B(n_484),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_645),
.A2(n_549),
.B(n_611),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_722),
.B(n_579),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_741),
.A2(n_514),
.B1(n_583),
.B2(n_614),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_657),
.A2(n_484),
.B1(n_602),
.B2(n_603),
.Y(n_792)
);

OAI321xp33_ASAP7_75t_L g793 ( 
.A1(n_653),
.A2(n_564),
.A3(n_568),
.B1(n_556),
.B2(n_544),
.C(n_603),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_631),
.B(n_602),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_754),
.B(n_608),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_674),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_630),
.A2(n_617),
.B(n_611),
.C(n_594),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_619),
.B(n_514),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_620),
.A2(n_621),
.B1(n_666),
.B2(n_685),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_677),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_595),
.C(n_594),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_654),
.B(n_633),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_704),
.B(n_579),
.Y(n_803)
);

BUFx5_ASAP7_75t_L g804 ( 
.A(n_751),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_518),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_688),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_639),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_690),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_766),
.A2(n_537),
.B(n_527),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_648),
.B(n_578),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_672),
.B(n_578),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_696),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_672),
.A2(n_527),
.B1(n_492),
.B2(n_609),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_684),
.A2(n_697),
.B(n_693),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_695),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_644),
.Y(n_817)
);

AOI21x1_ASAP7_75t_L g818 ( 
.A1(n_663),
.A2(n_609),
.B(n_242),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_755),
.B(n_50),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_684),
.A2(n_242),
.B(n_168),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_709),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_725),
.B(n_50),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_735),
.B(n_739),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_718),
.A2(n_52),
.B(n_242),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_693),
.A2(n_168),
.B(n_56),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_649),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_697),
.A2(n_98),
.B(n_57),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_630),
.A2(n_59),
.B(n_61),
.C(n_68),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_705),
.A2(n_70),
.B(n_75),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_625),
.A2(n_77),
.B(n_113),
.C(n_118),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_712),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_718),
.A2(n_121),
.B(n_131),
.C(n_133),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_713),
.B(n_149),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_686),
.A2(n_626),
.B(n_730),
.C(n_747),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_760),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_705),
.A2(n_729),
.B(n_720),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_706),
.A2(n_146),
.B(n_148),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_716),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_744),
.A2(n_762),
.B(n_764),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_716),
.A2(n_720),
.B(n_727),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_708),
.B(n_750),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_751),
.A2(n_722),
.B1(n_638),
.B2(n_703),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_741),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_765),
.B(n_636),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_698),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_L g846 ( 
.A1(n_623),
.A2(n_652),
.B(n_646),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_619),
.A2(n_622),
.B1(n_661),
.B2(n_642),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_724),
.A2(n_743),
.B(n_727),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_741),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_658),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_656),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_744),
.A2(n_731),
.B(n_635),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_683),
.A2(n_661),
.B(n_642),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_628),
.B(n_655),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_767),
.A2(n_757),
.B(n_745),
.C(n_748),
.Y(n_855)
);

BUFx4f_ASAP7_75t_L g856 ( 
.A(n_665),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_683),
.B(n_679),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_668),
.A2(n_717),
.B1(n_710),
.B2(n_719),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_656),
.Y(n_859)
);

AOI22x1_ASAP7_75t_L g860 ( 
.A1(n_658),
.A2(n_676),
.B1(n_679),
.B2(n_673),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_715),
.A2(n_734),
.B(n_733),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_721),
.A2(n_732),
.B(n_728),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_655),
.B(n_665),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_664),
.B(n_680),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_651),
.A2(n_701),
.B(n_667),
.C(n_699),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_671),
.A2(n_675),
.B(n_746),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_658),
.A2(n_682),
.B(n_761),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_761),
.A2(n_738),
.B(n_742),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_691),
.A2(n_692),
.B(n_694),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_689),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_740),
.A2(n_624),
.B(n_752),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_737),
.B(n_749),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_726),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_753),
.B(n_758),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_698),
.A2(n_759),
.B1(n_723),
.B2(n_740),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_723),
.B(n_678),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_756),
.A2(n_637),
.B(n_632),
.C(n_700),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_637),
.A2(n_645),
.B(n_643),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_714),
.B(n_485),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_704),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_660),
.A2(n_707),
.B(n_662),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_660),
.A2(n_707),
.B(n_662),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_660),
.A2(n_707),
.B(n_662),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_637),
.A2(n_632),
.B(n_700),
.C(n_643),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_687),
.B(n_643),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_714),
.B(n_485),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_695),
.Y(n_889)
);

AND2x2_ASAP7_75t_SL g890 ( 
.A(n_751),
.B(n_543),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_722),
.B(n_659),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_659),
.A2(n_663),
.B(n_662),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_641),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_618),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_637),
.A2(n_645),
.B(n_643),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_629),
.B(n_532),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_618),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_648),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_637),
.A2(n_632),
.B(n_700),
.C(n_643),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_629),
.B(n_335),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_637),
.A2(n_643),
.B1(n_687),
.B2(n_621),
.Y(n_901)
);

OAI321xp33_ASAP7_75t_L g902 ( 
.A1(n_711),
.A2(n_763),
.A3(n_653),
.B1(n_668),
.B2(n_637),
.C(n_670),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_687),
.B(n_643),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_641),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_637),
.A2(n_643),
.B1(n_687),
.B2(n_621),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_714),
.B(n_485),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_687),
.B(n_643),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_714),
.A2(n_736),
.B1(n_668),
.B2(n_711),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_629),
.B(n_335),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_711),
.A2(n_763),
.B(n_754),
.C(n_637),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_704),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_687),
.B(n_643),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_769),
.B(n_881),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_903),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_790),
.B(n_910),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_907),
.B(n_912),
.Y(n_916)
);

AO31x2_ASAP7_75t_L g917 ( 
.A1(n_787),
.A2(n_855),
.A3(n_785),
.B(n_905),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_802),
.A2(n_847),
.B1(n_821),
.B2(n_823),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_770),
.A2(n_899),
.B(n_886),
.C(n_834),
.Y(n_919)
);

AO21x1_ASAP7_75t_L g920 ( 
.A1(n_824),
.A2(n_879),
.B(n_883),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_890),
.B(n_864),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_882),
.B(n_911),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_888),
.B(n_906),
.Y(n_923)
);

OAI21x1_ASAP7_75t_SL g924 ( 
.A1(n_824),
.A2(n_905),
.B(n_901),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_795),
.A2(n_885),
.B(n_884),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_877),
.Y(n_926)
);

AOI21xp33_ASAP7_75t_L g927 ( 
.A1(n_858),
.A2(n_902),
.B(n_900),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_871),
.B(n_908),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_839),
.A2(n_852),
.B(n_777),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_839),
.A2(n_852),
.B(n_880),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_790),
.B(n_811),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_880),
.A2(n_895),
.B(n_789),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_790),
.B(n_771),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_902),
.A2(n_865),
.B(n_776),
.C(n_846),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_812),
.A2(n_842),
.B(n_858),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_790),
.B(n_783),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_SL g937 ( 
.A(n_909),
.B(n_779),
.C(n_801),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_768),
.B(n_774),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_877),
.B(n_856),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_778),
.A2(n_870),
.B(n_866),
.Y(n_941)
);

OAI22x1_ASAP7_75t_L g942 ( 
.A1(n_792),
.A2(n_798),
.B1(n_876),
.B2(n_819),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_796),
.B(n_800),
.Y(n_943)
);

OAI21x1_ASAP7_75t_SL g944 ( 
.A1(n_892),
.A2(n_797),
.B(n_895),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_868),
.A2(n_867),
.B(n_872),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_874),
.A2(n_772),
.B(n_828),
.C(n_842),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_806),
.B(n_807),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_808),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_804),
.B(n_794),
.Y(n_949)
);

AOI21xp33_ASAP7_75t_L g950 ( 
.A1(n_896),
.A2(n_772),
.B(n_873),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_815),
.A2(n_836),
.B(n_848),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_809),
.B(n_813),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_799),
.A2(n_832),
.B(n_830),
.C(n_784),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_840),
.A2(n_857),
.B(n_782),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_893),
.B(n_904),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_804),
.B(n_775),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_788),
.B(n_898),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_785),
.A2(n_799),
.B1(n_891),
.B2(n_835),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_875),
.B(n_891),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_805),
.B(n_819),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_863),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_817),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_793),
.A2(n_833),
.B(n_810),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_775),
.Y(n_964)
);

BUFx2_ASAP7_75t_SL g965 ( 
.A(n_845),
.Y(n_965)
);

BUFx2_ASAP7_75t_SL g966 ( 
.A(n_845),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_891),
.B(n_856),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_841),
.B(n_780),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_826),
.B(n_822),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_838),
.B(n_804),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_804),
.B(n_859),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_803),
.A2(n_814),
.B(n_850),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_SL g973 ( 
.A(n_889),
.B(n_878),
.C(n_831),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_851),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_816),
.B(n_843),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_825),
.A2(n_820),
.B(n_837),
.Y(n_976)
);

OAI33xp33_ASAP7_75t_L g977 ( 
.A1(n_894),
.A2(n_897),
.A3(n_844),
.B1(n_793),
.B2(n_849),
.B3(n_804),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_827),
.A2(n_829),
.B(n_869),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_877),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_850),
.B(n_869),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_887),
.B(n_903),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_860),
.A2(n_773),
.B(n_853),
.Y(n_982)
);

AO31x2_ASAP7_75t_L g983 ( 
.A1(n_787),
.A2(n_910),
.A3(n_855),
.B(n_785),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_887),
.B(n_903),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_887),
.B(n_903),
.Y(n_986)
);

OAI21x1_ASAP7_75t_SL g987 ( 
.A1(n_824),
.A2(n_886),
.B(n_770),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_802),
.A2(n_795),
.B(n_883),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_768),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_SL g991 ( 
.A1(n_824),
.A2(n_802),
.B(n_751),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_SL g994 ( 
.A1(n_824),
.A2(n_802),
.B(n_751),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_779),
.B(n_629),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_843),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_910),
.A2(n_770),
.B(n_899),
.C(n_886),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_910),
.A2(n_770),
.B(n_899),
.C(n_886),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_787),
.A2(n_818),
.B(n_777),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_889),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_887),
.B(n_903),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_802),
.A2(n_795),
.B(n_883),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_877),
.Y(n_1003)
);

AO31x2_ASAP7_75t_L g1004 ( 
.A1(n_787),
.A2(n_910),
.A3(n_855),
.B(n_785),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_889),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_889),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_887),
.B(n_903),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_802),
.A2(n_795),
.B(n_883),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_768),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_860),
.A2(n_839),
.B(n_852),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_790),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_887),
.B(n_903),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_845),
.B(n_498),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_SL g1015 ( 
.A1(n_802),
.A2(n_822),
.B(n_631),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_768),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_887),
.B(n_903),
.Y(n_1017)
);

NAND2x1_ASAP7_75t_L g1018 ( 
.A(n_869),
.B(n_877),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_910),
.A2(n_770),
.B(n_899),
.C(n_886),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_SL g1020 ( 
.A1(n_824),
.A2(n_802),
.B(n_751),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_853),
.A2(n_862),
.B(n_861),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_860),
.A2(n_839),
.B(n_852),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_824),
.A2(n_839),
.B(n_787),
.C(n_802),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_882),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_882),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_860),
.A2(n_839),
.B(n_852),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_769),
.B(n_485),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_889),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_887),
.B(n_903),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_768),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_887),
.B(n_903),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_781),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_860),
.A2(n_839),
.B(n_852),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_787),
.A2(n_910),
.A3(n_855),
.B(n_785),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_1000),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_996),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_957),
.B(n_913),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_984),
.A2(n_992),
.B(n_990),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1005),
.Y(n_1039)
);

HAxp5_ASAP7_75t_L g1040 ( 
.A(n_995),
.B(n_937),
.CON(n_1040),
.SN(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_1011),
.B(n_922),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_1024),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_914),
.B(n_916),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_940),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_981),
.B(n_985),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_927),
.A2(n_994),
.B(n_991),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1020),
.A2(n_1023),
.B(n_919),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_926),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_986),
.A2(n_1001),
.B1(n_1031),
.B2(n_1029),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_1024),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1007),
.A2(n_1013),
.B1(n_1017),
.B2(n_918),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1027),
.B(n_1006),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_960),
.B(n_923),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_958),
.A2(n_1019),
.B1(n_998),
.B2(n_997),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_967),
.B(n_965),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_993),
.A2(n_1021),
.B(n_1012),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_973),
.B(n_922),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1028),
.B(n_921),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_958),
.A2(n_997),
.B1(n_1019),
.B2(n_998),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_SL g1060 ( 
.A1(n_928),
.A2(n_924),
.B1(n_936),
.B2(n_915),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_919),
.A2(n_953),
.B(n_934),
.C(n_987),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_938),
.B(n_943),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_989),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_934),
.B(n_953),
.C(n_915),
.Y(n_1064)
);

OAI321xp33_ASAP7_75t_L g1065 ( 
.A1(n_946),
.A2(n_1002),
.A3(n_1008),
.B1(n_988),
.B2(n_925),
.C(n_941),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_922),
.Y(n_1066)
);

INVx6_ASAP7_75t_L g1067 ( 
.A(n_1025),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_926),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_947),
.B(n_952),
.Y(n_1069)
);

OA21x2_ASAP7_75t_L g1070 ( 
.A1(n_1010),
.A2(n_1033),
.B(n_1022),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1009),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_955),
.A2(n_946),
.B1(n_933),
.B2(n_1030),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_975),
.B(n_1025),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_959),
.B(n_935),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1016),
.B(n_950),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_974),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_969),
.A2(n_931),
.B1(n_961),
.B2(n_1014),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_996),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_942),
.B(n_968),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_926),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_961),
.A2(n_970),
.B1(n_971),
.B2(n_939),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_932),
.A2(n_930),
.B(n_1033),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_948),
.B(n_1032),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_948),
.Y(n_1084)
);

CKINVDCx16_ASAP7_75t_R g1085 ( 
.A(n_966),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_979),
.B(n_964),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_977),
.B(n_964),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_962),
.B(n_1032),
.Y(n_1088)
);

CKINVDCx6p67_ASAP7_75t_R g1089 ( 
.A(n_1003),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_956),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1003),
.B(n_1034),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1018),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_980),
.B1(n_930),
.B2(n_956),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_917),
.B(n_1034),
.Y(n_1094)
);

BUFx4f_ASAP7_75t_L g1095 ( 
.A(n_1015),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_983),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_949),
.B(n_972),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_980),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_983),
.B(n_1034),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_963),
.A2(n_944),
.B1(n_932),
.B2(n_929),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_917),
.B(n_983),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_963),
.A2(n_929),
.B1(n_1010),
.B2(n_1026),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_1034),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_983),
.B(n_1004),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_954),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_1004),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1004),
.B(n_917),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1004),
.B(n_917),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_951),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_945),
.B(n_999),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_982),
.A2(n_927),
.B(n_598),
.C(n_802),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_978),
.B(n_976),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_976),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1011),
.B(n_967),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_940),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1000),
.Y(n_1116)
);

INVxp67_ASAP7_75t_SL g1117 ( 
.A(n_914),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_1024),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1011),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_940),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_1024),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_996),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1011),
.B(n_979),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1011),
.B(n_922),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_984),
.A2(n_992),
.B(n_990),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1000),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_940),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_995),
.A2(n_783),
.B1(n_927),
.B2(n_580),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_996),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_SL g1130 ( 
.A(n_1011),
.B(n_926),
.Y(n_1130)
);

OAI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_927),
.A2(n_598),
.B(n_580),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_933),
.B(n_914),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_984),
.A2(n_992),
.B(n_990),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_957),
.B(n_913),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_1024),
.B(n_704),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_984),
.A2(n_992),
.B(n_990),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_920),
.A2(n_927),
.B(n_824),
.C(n_1023),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1011),
.B(n_979),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1011),
.B(n_922),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_914),
.A2(n_637),
.B1(n_910),
.B2(n_916),
.Y(n_1140)
);

CKINVDCx8_ASAP7_75t_R g1141 ( 
.A(n_965),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1011),
.B(n_922),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_995),
.B(n_629),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_926),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_1000),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1011),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_927),
.A2(n_598),
.B(n_802),
.C(n_937),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_926),
.Y(n_1148)
);

AOI221x1_ASAP7_75t_L g1149 ( 
.A1(n_927),
.A2(n_934),
.B1(n_910),
.B2(n_946),
.C(n_824),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_995),
.B(n_629),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_914),
.B(n_916),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_914),
.A2(n_637),
.B1(n_910),
.B2(n_916),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_984),
.A2(n_992),
.B(n_990),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_940),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_995),
.B(n_629),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_914),
.A2(n_637),
.B1(n_910),
.B2(n_916),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1145),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1099),
.B(n_1104),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1067),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1038),
.A2(n_1125),
.B(n_1056),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1063),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1117),
.B(n_1043),
.Y(n_1162)
);

AO21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1047),
.A2(n_1046),
.B(n_1094),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1071),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1115),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1120),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1109),
.A2(n_1054),
.B1(n_1059),
.B2(n_1064),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1127),
.Y(n_1168)
);

BUFx2_ASAP7_75t_R g1169 ( 
.A(n_1036),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1108),
.B(n_1107),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1068),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1107),
.B(n_1105),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1043),
.B(n_1151),
.Y(n_1173)
);

CKINVDCx8_ASAP7_75t_R g1174 ( 
.A(n_1085),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_1054),
.A2(n_1059),
.B(n_1061),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1131),
.A2(n_1128),
.B1(n_1064),
.B2(n_1079),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1097),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1067),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_1129),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1151),
.B(n_1049),
.Y(n_1180)
);

INVx8_ASAP7_75t_L g1181 ( 
.A(n_1080),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1049),
.A2(n_1051),
.B1(n_1075),
.B2(n_1150),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_1122),
.Y(n_1183)
);

AOI222xp33_ASAP7_75t_L g1184 ( 
.A1(n_1051),
.A2(n_1045),
.B1(n_1156),
.B2(n_1140),
.C1(n_1152),
.C2(n_1134),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1047),
.B(n_1106),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1154),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1039),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1147),
.A2(n_1060),
.B1(n_1156),
.B2(n_1152),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1075),
.A2(n_1155),
.B1(n_1143),
.B2(n_1058),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1097),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1035),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1076),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1140),
.A2(n_1072),
.B1(n_1087),
.B2(n_1062),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1037),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1116),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1133),
.A2(n_1153),
.B(n_1136),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1072),
.A2(n_1087),
.B1(n_1069),
.B2(n_1077),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1149),
.A2(n_1111),
.B(n_1130),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1096),
.B(n_1091),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1084),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1042),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1126),
.B(n_1052),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1124),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1132),
.B(n_1053),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1068),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1083),
.Y(n_1206)
);

CKINVDCx14_ASAP7_75t_R g1207 ( 
.A(n_1073),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1074),
.B(n_1101),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1097),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1088),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1082),
.A2(n_1065),
.B(n_1137),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1118),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1066),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1078),
.A2(n_1098),
.B1(n_1057),
.B2(n_1065),
.Y(n_1214)
);

CKINVDCx6p67_ASAP7_75t_R g1215 ( 
.A(n_1055),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1141),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1114),
.B(n_1074),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1086),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1102),
.A2(n_1100),
.B(n_1110),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1077),
.A2(n_1101),
.B1(n_1094),
.B2(n_1103),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_1050),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_SL g1222 ( 
.A(n_1121),
.Y(n_1222)
);

AOI22x1_ASAP7_75t_SL g1223 ( 
.A1(n_1040),
.A2(n_1119),
.B1(n_1146),
.B2(n_1092),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1070),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1095),
.A2(n_1081),
.B(n_1093),
.Y(n_1225)
);

BUFx2_ASAP7_75t_R g1226 ( 
.A(n_1048),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1144),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1093),
.B(n_1081),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_1112),
.A2(n_1138),
.B(n_1123),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1144),
.Y(n_1230)
);

AO21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1095),
.A2(n_1113),
.B(n_1112),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1148),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1148),
.Y(n_1233)
);

BUFx2_ASAP7_75t_SL g1234 ( 
.A(n_1139),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1148),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1142),
.A2(n_1135),
.B1(n_1138),
.B2(n_1123),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1048),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1089),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1113),
.A2(n_927),
.B1(n_890),
.B2(n_772),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1067),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1090),
.B(n_1041),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1044),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1044),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1054),
.A2(n_783),
.B1(n_927),
.B2(n_792),
.Y(n_1244)
);

BUFx2_ASAP7_75t_R g1245 ( 
.A(n_1036),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1145),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1131),
.A2(n_927),
.B1(n_890),
.B2(n_772),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1145),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1109),
.A2(n_791),
.B1(n_513),
.B2(n_474),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1090),
.B(n_1041),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1067),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_SL g1253 ( 
.A(n_1129),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1117),
.B(n_1043),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1062),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1044),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1224),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1177),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1208),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1187),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1208),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1217),
.B(n_1229),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1190),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1175),
.A2(n_1160),
.B(n_1188),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1200),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1158),
.B(n_1185),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1206),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1209),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1158),
.B(n_1185),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1183),
.Y(n_1270)
);

BUFx8_ASAP7_75t_L g1271 ( 
.A(n_1249),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1228),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1163),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1228),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1256),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1215),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1174),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1180),
.B(n_1255),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1209),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1161),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1215),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1213),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_SL g1285 ( 
.A(n_1249),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1231),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1164),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1244),
.A2(n_1225),
.B(n_1229),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1199),
.B(n_1165),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1196),
.A2(n_1160),
.B(n_1211),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1199),
.B(n_1166),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1198),
.A2(n_1162),
.B(n_1254),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1218),
.B(n_1194),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1168),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1167),
.A2(n_1193),
.B(n_1197),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1186),
.B(n_1242),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1198),
.A2(n_1192),
.B(n_1247),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1195),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1218),
.B(n_1217),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1243),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1253),
.B(n_1221),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1191),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1211),
.A2(n_1219),
.B(n_1176),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1210),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1219),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1219),
.A2(n_1239),
.B(n_1175),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1227),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1220),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1189),
.B(n_1173),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1237),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1237),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1214),
.A2(n_1235),
.B(n_1232),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1207),
.B(n_1204),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1207),
.B(n_1241),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1233),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1266),
.B(n_1171),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1297),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1290),
.A2(n_1248),
.B(n_1236),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1278),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1297),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1280),
.B(n_1201),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1297),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1286),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1257),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1265),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1258),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1276),
.B(n_1202),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1265),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1277),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1277),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1303),
.A2(n_1212),
.B1(n_1157),
.B2(n_1246),
.C(n_1159),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1258),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1306),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1295),
.B(n_1223),
.C(n_1250),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1276),
.B(n_1252),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1263),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1266),
.B(n_1205),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1269),
.B(n_1205),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1269),
.B(n_1205),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1303),
.A2(n_1174),
.B1(n_1221),
.B2(n_1226),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1259),
.B(n_1230),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1278),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1264),
.A2(n_1238),
.B(n_1251),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1286),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1274),
.B(n_1252),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1263),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1275),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1289),
.B(n_1230),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1306),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1289),
.B(n_1230),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1291),
.B(n_1240),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1283),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1283),
.Y(n_1356)
);

AOI222xp33_ASAP7_75t_L g1357 ( 
.A1(n_1309),
.A2(n_1157),
.B1(n_1246),
.B2(n_1222),
.C1(n_1183),
.C2(n_1251),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1286),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1264),
.A2(n_1159),
.B1(n_1178),
.B2(n_1234),
.C(n_1203),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1345),
.B(n_1272),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1320),
.B(n_1283),
.Y(n_1361)
);

NAND4xp25_ASAP7_75t_L g1362 ( 
.A(n_1335),
.B(n_1309),
.C(n_1301),
.D(n_1275),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1345),
.B(n_1272),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1335),
.B(n_1308),
.C(n_1316),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1328),
.B(n_1260),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1328),
.B(n_1298),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1345),
.B(n_1273),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1341),
.A2(n_1314),
.B1(n_1282),
.B2(n_1300),
.C(n_1294),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1336),
.B(n_1292),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1325),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1317),
.B(n_1273),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1341),
.A2(n_1357),
.B(n_1332),
.Y(n_1372)
);

OAI221xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1332),
.A2(n_1293),
.B1(n_1314),
.B2(n_1262),
.C(n_1310),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1322),
.B(n_1292),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1344),
.B(n_1284),
.C(n_1302),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1344),
.B(n_1311),
.C(n_1312),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1357),
.B(n_1311),
.C(n_1312),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1338),
.B(n_1339),
.Y(n_1378)
);

AOI21xp33_ASAP7_75t_L g1379 ( 
.A1(n_1346),
.A2(n_1288),
.B(n_1313),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1359),
.A2(n_1315),
.B(n_1279),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1334),
.A2(n_1307),
.B(n_1304),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1351),
.B(n_1296),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1359),
.A2(n_1315),
.B(n_1279),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1353),
.B(n_1296),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1327),
.B(n_1268),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1339),
.B(n_1268),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1348),
.B(n_1300),
.C(n_1287),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1319),
.A2(n_1288),
.B1(n_1307),
.B2(n_1313),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1287),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1340),
.B(n_1294),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_L g1391 ( 
.A(n_1348),
.B(n_1267),
.C(n_1305),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1340),
.B(n_1267),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1346),
.A2(n_1288),
.B1(n_1307),
.B2(n_1321),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1318),
.A2(n_1262),
.B1(n_1306),
.B2(n_1299),
.C(n_1288),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1327),
.B(n_1281),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1368),
.B(n_1333),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1372),
.B(n_1354),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1370),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1378),
.B(n_1334),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1378),
.B(n_1352),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1387),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1371),
.B(n_1352),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1371),
.B(n_1346),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1387),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1360),
.B(n_1346),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1369),
.B(n_1326),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1391),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1360),
.B(n_1342),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1391),
.Y(n_1409)
);

AND2x4_ASAP7_75t_SL g1410 ( 
.A(n_1363),
.B(n_1324),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1385),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1375),
.B(n_1326),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1375),
.B(n_1329),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1365),
.B(n_1337),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1389),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1367),
.B(n_1329),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1376),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1390),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1386),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1385),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1392),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_SL g1422 ( 
.A(n_1361),
.B(n_1347),
.Y(n_1422)
);

NAND2x1_ASAP7_75t_L g1423 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1366),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1374),
.B(n_1330),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1416),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1416),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1397),
.B(n_1372),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1401),
.B(n_1382),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1405),
.B(n_1337),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1405),
.B(n_1349),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1401),
.B(n_1384),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1403),
.B(n_1350),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1398),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1410),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1403),
.B(n_1350),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1412),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1412),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1413),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1403),
.B(n_1395),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1397),
.A2(n_1362),
.B1(n_1381),
.B2(n_1379),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1398),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1399),
.B(n_1364),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1423),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1413),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1417),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1404),
.B(n_1330),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1404),
.B(n_1331),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1425),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1425),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1407),
.B(n_1394),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1399),
.B(n_1400),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1398),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1415),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1417),
.A2(n_1321),
.B1(n_1323),
.B2(n_1377),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1415),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1407),
.B(n_1331),
.Y(n_1457)
);

AND2x6_ASAP7_75t_SL g1458 ( 
.A(n_1409),
.B(n_1271),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1418),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1428),
.A2(n_1396),
.B(n_1409),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1428),
.B(n_1424),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1437),
.B(n_1424),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1444),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1438),
.B(n_1396),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1406),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1439),
.B(n_1418),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1458),
.B(n_1285),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1454),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1421),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1458),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1445),
.B(n_1421),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1452),
.B(n_1419),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1452),
.B(n_1419),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1434),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1429),
.B(n_1271),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1441),
.A2(n_1362),
.B1(n_1393),
.B2(n_1381),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1454),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1434),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1445),
.B(n_1420),
.Y(n_1486)
);

NAND4xp25_ASAP7_75t_L g1487 ( 
.A(n_1441),
.B(n_1377),
.C(n_1414),
.D(n_1411),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1452),
.B(n_1419),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1434),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1410),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1442),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1432),
.B(n_1406),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1444),
.Y(n_1494)
);

OR2x6_ASAP7_75t_SL g1495 ( 
.A(n_1451),
.B(n_1446),
.Y(n_1495)
);

OAI21xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1451),
.A2(n_1400),
.B(n_1402),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1433),
.B(n_1419),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1455),
.A2(n_1388),
.B1(n_1383),
.B2(n_1380),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1447),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1429),
.B(n_1271),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1435),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1456),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1465),
.B(n_1440),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1482),
.A2(n_1455),
.B1(n_1446),
.B2(n_1459),
.C(n_1373),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1473),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1483),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1483),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1462),
.B(n_1446),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1495),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1470),
.B(n_1446),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1470),
.B(n_1459),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1501),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1271),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1465),
.B(n_1440),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1501),
.B(n_1459),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1495),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1493),
.B(n_1459),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_L g1520 ( 
.A(n_1475),
.B(n_1179),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1503),
.Y(n_1522)
);

INVx5_ASAP7_75t_L g1523 ( 
.A(n_1466),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1472),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1482),
.B(n_1498),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1503),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1464),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1467),
.B(n_1433),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1468),
.B(n_1436),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1468),
.B(n_1436),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1463),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1492),
.B(n_1426),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1534)
);

AOI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1487),
.A2(n_1449),
.B1(n_1450),
.B2(n_1457),
.C(n_1448),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1461),
.A2(n_1453),
.B(n_1442),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1466),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1426),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_R g1539 ( 
.A(n_1494),
.B(n_1216),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_L g1540 ( 
.A(n_1525),
.B(n_1498),
.C(n_1496),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1505),
.A2(n_1496),
.B1(n_1469),
.B2(n_1499),
.C(n_1450),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1532),
.B(n_1502),
.Y(n_1542)
);

OAI32xp33_ASAP7_75t_L g1543 ( 
.A1(n_1511),
.A2(n_1484),
.A3(n_1466),
.B1(n_1486),
.B2(n_1500),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1536),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1518),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1534),
.B(n_1471),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1477),
.Y(n_1547)
);

OAI322xp33_ASAP7_75t_L g1548 ( 
.A1(n_1518),
.A2(n_1476),
.A3(n_1474),
.B1(n_1484),
.B2(n_1448),
.C1(n_1447),
.C2(n_1457),
.Y(n_1548)
);

XNOR2x1_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1536),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1514),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1536),
.A2(n_1380),
.B1(n_1383),
.B2(n_1491),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1508),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1524),
.B(n_1270),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1536),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1509),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1510),
.A2(n_1485),
.B(n_1479),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1510),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1509),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1533),
.A2(n_1484),
.B(n_1494),
.C(n_1481),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1522),
.Y(n_1563)
);

AOI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1512),
.A2(n_1485),
.B(n_1479),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1169),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1556),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1556),
.A2(n_1535),
.B1(n_1489),
.B2(n_1491),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1545),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1540),
.A2(n_1504),
.B1(n_1521),
.B2(n_1516),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1554),
.B(n_1516),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1553),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1562),
.B(n_1521),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1549),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1559),
.B(n_1527),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1557),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1565),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_SL g1581 ( 
.A(n_1543),
.B(n_1539),
.C(n_1537),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1546),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1550),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1551),
.A2(n_1534),
.B1(n_1512),
.B2(n_1513),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_L g1586 ( 
.A(n_1576),
.B(n_1541),
.C(n_1559),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1569),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1567),
.A2(n_1564),
.B1(n_1558),
.B2(n_1561),
.C(n_1513),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1585),
.A2(n_1548),
.B(n_1542),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1570),
.A2(n_1547),
.B(n_1507),
.Y(n_1590)
);

AOI21xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1577),
.A2(n_1563),
.B(n_1560),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1581),
.B(n_1523),
.C(n_1517),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1517),
.B(n_1519),
.C(n_1522),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1580),
.B(n_1519),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1568),
.A2(n_1517),
.B1(n_1489),
.B2(n_1526),
.Y(n_1595)
);

NOR4xp25_ASAP7_75t_L g1596 ( 
.A(n_1582),
.B(n_1526),
.C(n_1506),
.D(n_1528),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1583),
.B(n_1523),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1575),
.Y(n_1598)
);

NOR4xp25_ASAP7_75t_L g1599 ( 
.A(n_1593),
.B(n_1582),
.C(n_1566),
.D(n_1584),
.Y(n_1599)
);

OAI211xp5_ASAP7_75t_L g1600 ( 
.A1(n_1596),
.A2(n_1566),
.B(n_1572),
.C(n_1578),
.Y(n_1600)
);

OAI211xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1589),
.A2(n_1571),
.B(n_1584),
.C(n_1583),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1597),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1586),
.B(n_1574),
.C(n_1573),
.Y(n_1603)
);

NAND5xp2_ASAP7_75t_L g1604 ( 
.A(n_1594),
.B(n_1575),
.C(n_1579),
.D(n_1528),
.E(n_1531),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1591),
.B(n_1530),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1592),
.B(n_1481),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1590),
.B(n_1530),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1588),
.B(n_1523),
.C(n_1531),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1601),
.A2(n_1595),
.B1(n_1538),
.B2(n_1523),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1598),
.Y(n_1610)
);

NOR3xp33_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1216),
.C(n_1538),
.Y(n_1611)
);

OA22x2_ASAP7_75t_L g1612 ( 
.A1(n_1602),
.A2(n_1481),
.B1(n_1490),
.B2(n_1435),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1604),
.B(n_1490),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1610),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1611),
.A2(n_1599),
.B1(n_1608),
.B2(n_1600),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1612),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1613),
.B(n_1605),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1609),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1612),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1616),
.B(n_1619),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1614),
.B(n_1606),
.Y(n_1621)
);

NOR3xp33_ASAP7_75t_L g1622 ( 
.A(n_1617),
.B(n_1607),
.C(n_1245),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_L g1623 ( 
.A(n_1618),
.B(n_1178),
.C(n_1442),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1615),
.B(n_1478),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1621),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1620),
.Y(n_1626)
);

NAND3x1_ASAP7_75t_L g1627 ( 
.A(n_1622),
.B(n_1488),
.C(n_1478),
.Y(n_1627)
);

OA22x2_ASAP7_75t_L g1628 ( 
.A1(n_1625),
.A2(n_1624),
.B1(n_1623),
.B2(n_1490),
.Y(n_1628)
);

NOR4xp25_ASAP7_75t_L g1629 ( 
.A(n_1628),
.B(n_1626),
.C(n_1627),
.D(n_1449),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1629),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1629),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1630),
.A2(n_1427),
.B1(n_1488),
.B2(n_1497),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1631),
.A2(n_1460),
.B(n_1456),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1633),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1632),
.B(n_1497),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1634),
.B(n_1453),
.C(n_1460),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1636),
.A2(n_1635),
.B1(n_1435),
.B2(n_1431),
.Y(n_1637)
);

OAI221xp5_ASAP7_75t_R g1638 ( 
.A1(n_1637),
.A2(n_1181),
.B1(n_1422),
.B2(n_1427),
.C(n_1430),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1638),
.A2(n_1355),
.B(n_1356),
.C(n_1343),
.Y(n_1639)
);


endmodule