module fake_ibex_12_n_1059 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1059);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1059;

wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1031;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_1018;
wire n_1044;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_283;
wire n_366;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_899;
wire n_843;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_807;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_890;
wire n_921;
wire n_912;
wire n_874;
wire n_1058;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_984;
wire n_1000;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g198 ( 
.A(n_39),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_58),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_9),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_47),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_56),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_46),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_35),
.B(n_69),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_79),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_157),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_123),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_124),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_46),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_110),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_172),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_60),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_34),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_140),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_119),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_54),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_26),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_32),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_32),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_121),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_41),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_161),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_43),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_77),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_67),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_131),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_17),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_106),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_114),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_104),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_78),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_111),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_175),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_91),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_156),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_126),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_152),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_169),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_163),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_21),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_185),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_99),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_83),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_48),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_75),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_45),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_134),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_160),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_45),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_130),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_117),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_166),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_48),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_147),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_87),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_133),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_11),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_74),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_158),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_146),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_109),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_165),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_93),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_6),
.Y(n_316)
);

INVx4_ASAP7_75t_R g317 ( 
.A(n_81),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_30),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_60),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_144),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_193),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_112),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_190),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_37),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_120),
.B(n_186),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_11),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_164),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_96),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_95),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_4),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_30),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_137),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_155),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_238),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_203),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_1),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_217),
.A2(n_68),
.B(n_66),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_213),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_216),
.B(n_3),
.Y(n_347)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_217),
.A2(n_71),
.B(n_70),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_216),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_242),
.B(n_4),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_213),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_205),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_226),
.A2(n_97),
.B(n_197),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_204),
.B(n_7),
.Y(n_356)
);

OR2x6_ASAP7_75t_L g357 ( 
.A(n_242),
.B(n_7),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_200),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_244),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_213),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_238),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_8),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_237),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_290),
.Y(n_369)
);

BUFx8_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_268),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_290),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_281),
.B(n_12),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_226),
.A2(n_101),
.B(n_195),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_213),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_220),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_281),
.B(n_14),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_228),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_228),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_208),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_228),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_275),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_212),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_214),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_219),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_285),
.B(n_15),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_228),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_200),
.B(n_72),
.Y(n_391)
);

NOR2x1_ASAP7_75t_L g392 ( 
.A(n_218),
.B(n_15),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_243),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_209),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_222),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_258),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_338),
.B(n_314),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_236),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_223),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_220),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_220),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_233),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_236),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_234),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_243),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_243),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_235),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_316),
.B(n_18),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_291),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_291),
.B(n_73),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_316),
.B(n_19),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_210),
.B(n_20),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_237),
.A2(n_319),
.B1(n_318),
.B2(n_201),
.Y(n_416)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_275),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_239),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_202),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_243),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_198),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

BUFx6f_ASAP7_75t_SL g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_395),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_353),
.B(n_253),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_313),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_389),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_355),
.B(n_276),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_362),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_399),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_232),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_419),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_370),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_240),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_368),
.A2(n_304),
.B1(n_207),
.B2(n_227),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_346),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_397),
.B(n_246),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_369),
.B(n_341),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_389),
.B(n_224),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_215),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_346),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_412),
.A2(n_241),
.B1(n_251),
.B2(n_249),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_412),
.B(n_247),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_385),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_370),
.B(n_254),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_370),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_416),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_369),
.B(n_259),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_341),
.B(n_252),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_344),
.B(n_256),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_417),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_351),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_260),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_340),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_375),
.B(n_279),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_391),
.B(n_379),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_357),
.B(n_265),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_394),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_354),
.A2(n_263),
.B(n_261),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_352),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g480 ( 
.A1(n_357),
.A2(n_304),
.B1(n_272),
.B2(n_283),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_398),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_352),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_363),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_360),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_366),
.B(n_269),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_L g486 ( 
.A1(n_357),
.A2(n_284),
.B1(n_286),
.B2(n_266),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_413),
.B(n_230),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_372),
.B(n_271),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_356),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_383),
.B(n_273),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_383),
.B(n_274),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_398),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_360),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_386),
.A2(n_296),
.B(n_289),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_360),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_386),
.B(n_277),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_345),
.B(n_230),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_345),
.B(n_230),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_387),
.B(n_294),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_387),
.B(n_295),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_410),
.B(n_320),
.C(n_307),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g504 ( 
.A1(n_354),
.A2(n_298),
.B(n_297),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_388),
.B(n_328),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_377),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_377),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_380),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_396),
.A2(n_401),
.B1(n_406),
.B2(n_404),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_411),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_380),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_391),
.B(n_312),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_380),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_326),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_382),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_382),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_349),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_404),
.B(n_299),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_382),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_365),
.Y(n_528)
);

AND2x2_ASAP7_75t_SL g529 ( 
.A(n_345),
.B(n_230),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_365),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_406),
.B(n_301),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_384),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_409),
.B(n_303),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_211),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_384),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_418),
.B(n_306),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_418),
.B(n_309),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_392),
.B(n_221),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_489),
.B(n_442),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_445),
.B(n_225),
.Y(n_540)
);

OAI221xp5_ASAP7_75t_L g541 ( 
.A1(n_494),
.A2(n_359),
.B1(n_421),
.B2(n_336),
.C(n_335),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_231),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_456),
.A2(n_278),
.B1(n_224),
.B2(n_229),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_465),
.B(n_392),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_444),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_486),
.A2(n_229),
.B1(n_248),
.B2(n_315),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_250),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_495),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_456),
.A2(n_315),
.B1(n_278),
.B2(n_300),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_498),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_468),
.B(n_311),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_255),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_446),
.B(n_450),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_463),
.B(n_264),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_471),
.B(n_339),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_469),
.B(n_378),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_503),
.B(n_324),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_475),
.A2(n_480),
.B1(n_486),
.B2(n_512),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_443),
.B(n_334),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_473),
.B(n_267),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_438),
.B(n_270),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_433),
.B(n_257),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_475),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_437),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_453),
.B(n_280),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_424),
.B(n_282),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_327),
.C(n_245),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_424),
.B(n_287),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_453),
.B(n_288),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_453),
.B(n_293),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_425),
.B(n_248),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_425),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_471),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_514),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_460),
.B(n_378),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_466),
.B(n_305),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_437),
.B(n_348),
.C(n_345),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_487),
.A2(n_300),
.B1(n_292),
.B2(n_257),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_451),
.B(n_308),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_480),
.B(n_310),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_462),
.B(n_321),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_479),
.B(n_257),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_518),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_457),
.B(n_332),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_436),
.B(n_333),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_518),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_462),
.B(n_337),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_519),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_447),
.B(n_330),
.C(n_403),
.Y(n_596)
);

NOR3x1_ASAP7_75t_L g597 ( 
.A(n_464),
.B(n_24),
.C(n_26),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_481),
.B(n_292),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_470),
.B(n_348),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_422),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_434),
.B(n_348),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_467),
.B(n_292),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_441),
.B(n_376),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_448),
.B(n_376),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_458),
.A2(n_402),
.B1(n_403),
.B2(n_323),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_528),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_530),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_458),
.A2(n_323),
.B1(n_408),
.B2(n_407),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_452),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_452),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_459),
.B(n_27),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_476),
.B(n_384),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_459),
.B(n_27),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

AND3x1_ASAP7_75t_L g617 ( 
.A(n_491),
.B(n_317),
.C(n_29),
.Y(n_617)
);

AOI22x1_ASAP7_75t_L g618 ( 
.A1(n_423),
.A2(n_420),
.B1(n_408),
.B2(n_407),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_511),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_513),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_497),
.B(n_390),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_538),
.B(n_390),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_526),
.B(n_390),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_492),
.A2(n_420),
.B1(n_408),
.B2(n_407),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_526),
.B(n_390),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_537),
.B(n_393),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_393),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_525),
.B(n_439),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_L g631 ( 
.A(n_488),
.B(n_28),
.C(n_29),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_488),
.B(n_407),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_539),
.B(n_490),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_602),
.A2(n_516),
.B(n_500),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_561),
.A2(n_536),
.B1(n_502),
.B2(n_533),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_561),
.A2(n_568),
.B1(n_546),
.B2(n_550),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_501),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_568),
.A2(n_502),
.B1(n_533),
.B2(n_501),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_543),
.A2(n_531),
.B1(n_500),
.B2(n_529),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_531),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_604),
.A2(n_516),
.B(n_499),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_563),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_595),
.B(n_499),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_606),
.A2(n_529),
.B(n_429),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_563),
.B(n_427),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_582),
.A2(n_504),
.B(n_477),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_600),
.A2(n_431),
.B(n_430),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_541),
.B(n_432),
.C(n_431),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_571),
.B(n_435),
.C(n_432),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_567),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_567),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_555),
.B(n_435),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_440),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_578),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_586),
.A2(n_535),
.B1(n_455),
.B2(n_527),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_593),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_599),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_552),
.A2(n_496),
.B1(n_523),
.B2(n_522),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_544),
.A2(n_496),
.B(n_523),
.C(n_522),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_584),
.A2(n_493),
.B1(n_521),
.B2(n_520),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_611),
.B(n_31),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_611),
.B(n_33),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_562),
.B(n_33),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_562),
.B(n_542),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_605),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_566),
.B(n_36),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_598),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_612),
.B(n_38),
.Y(n_671)
);

NAND2x1p5_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_38),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_599),
.B(n_42),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_560),
.A2(n_508),
.B(n_478),
.C(n_515),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_565),
.B(n_43),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_SL g676 ( 
.A(n_571),
.B(n_596),
.C(n_631),
.Y(n_676)
);

INVxp33_ASAP7_75t_SL g677 ( 
.A(n_581),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_588),
.B(n_44),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_608),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

NOR2x1_ASAP7_75t_L g681 ( 
.A(n_558),
.B(n_509),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_596),
.B(n_510),
.C(n_509),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_590),
.B(n_44),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_47),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_624),
.A2(n_510),
.B(n_532),
.C(n_517),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_580),
.B(n_49),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_630),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_630),
.B(n_49),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_603),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_624),
.A2(n_532),
.B(n_517),
.C(n_484),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_573),
.B(n_50),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_621),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_547),
.B(n_50),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_616),
.A2(n_482),
.B1(n_449),
.B2(n_53),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_569),
.B(n_574),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_621),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_620),
.B(n_51),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_628),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_631),
.A2(n_52),
.B(n_54),
.C(n_57),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_619),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_627),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_554),
.A2(n_135),
.B(n_192),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_621),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_558),
.B(n_59),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_613),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_564),
.B(n_61),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_558),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_587),
.A2(n_139),
.B(n_189),
.C(n_76),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_579),
.Y(n_710)
);

BUFx8_ASAP7_75t_L g711 ( 
.A(n_615),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_594),
.B(n_184),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_591),
.A2(n_80),
.B(n_82),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_585),
.A2(n_85),
.B(n_86),
.C(n_88),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_603),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_105),
.B(n_107),
.C(n_108),
.Y(n_716)
);

BUFx12f_ASAP7_75t_L g717 ( 
.A(n_597),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_583),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_540),
.B(n_127),
.Y(n_719)
);

BUFx8_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_557),
.B(n_129),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_548),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_592),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_622),
.A2(n_629),
.B(n_626),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_559),
.B(n_182),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_136),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_607),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_610),
.A3(n_623),
.B(n_614),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_720),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_720),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_650),
.B(n_632),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_651),
.B(n_572),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_644),
.A2(n_625),
.B(n_570),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_618),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_636),
.B(n_168),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_636),
.B(n_171),
.Y(n_737)
);

AND2x2_ASAP7_75t_SL g738 ( 
.A(n_687),
.B(n_174),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_653),
.B(n_176),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_658),
.B(n_179),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_639),
.A2(n_635),
.B1(n_708),
.B2(n_695),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_647),
.A2(n_637),
.B(n_633),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_670),
.B(n_640),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_668),
.B(n_705),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_639),
.A2(n_685),
.A3(n_661),
.B(n_728),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_694),
.B(n_649),
.C(n_675),
.Y(n_746)
);

CKINVDCx11_ASAP7_75t_R g747 ( 
.A(n_717),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_711),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_688),
.B(n_672),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_648),
.B(n_667),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_724),
.A2(n_638),
.B(n_643),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_679),
.B(n_680),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_655),
.B(n_678),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_711),
.B(n_681),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_654),
.Y(n_755)
);

AO31x2_ASAP7_75t_L g756 ( 
.A1(n_694),
.A2(n_674),
.A3(n_716),
.B(n_698),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_SL g757 ( 
.A1(n_708),
.A2(n_699),
.B(n_701),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_665),
.B(n_663),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_664),
.B(n_671),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_691),
.A2(n_683),
.B(n_684),
.C(n_693),
.Y(n_760)
);

BUFx10_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_682),
.A2(n_702),
.B(n_713),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_700),
.B(n_706),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_722),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_697),
.A2(n_669),
.B1(n_673),
.B2(n_715),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_659),
.B(n_692),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_707),
.A2(n_723),
.B1(n_718),
.B2(n_710),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_719),
.A2(n_721),
.B1(n_660),
.B2(n_673),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_712),
.B(n_722),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_659),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_727),
.B(n_725),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_727),
.B(n_703),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_692),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_714),
.B(n_709),
.C(n_662),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_656),
.A3(n_696),
.B(n_703),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_696),
.B(n_539),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_657),
.B(n_539),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_658),
.B(n_601),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_657),
.B(n_539),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_654),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_720),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_666),
.B(n_539),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_650),
.B(n_545),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_666),
.B(n_539),
.Y(n_785)
);

OA22x2_ASAP7_75t_L g786 ( 
.A1(n_636),
.A2(n_546),
.B1(n_398),
.B2(n_545),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_642),
.B(n_545),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_646),
.A2(n_504),
.B(n_477),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_720),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_644),
.A2(n_641),
.B(n_634),
.Y(n_790)
);

AOI21x1_ASAP7_75t_L g791 ( 
.A1(n_646),
.A2(n_504),
.B(n_477),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_690),
.A2(n_600),
.A3(n_644),
.B(n_641),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_652),
.B(n_567),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_642),
.B(n_545),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_720),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_SL g796 ( 
.A1(n_636),
.A2(n_561),
.B(n_708),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_634),
.A2(n_474),
.B(n_437),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_720),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_642),
.B(n_545),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_720),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_545),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_654),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_634),
.A2(n_474),
.B(n_437),
.Y(n_803)
);

AOI221xp5_ASAP7_75t_L g804 ( 
.A1(n_636),
.A2(n_561),
.B1(n_447),
.B2(n_541),
.C(n_571),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_636),
.A2(n_639),
.B1(n_456),
.B2(n_652),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_650),
.B(n_545),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_644),
.A2(n_641),
.B(n_634),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_720),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_690),
.A2(n_600),
.A3(n_644),
.B(n_641),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_666),
.B(n_539),
.Y(n_810)
);

AO31x2_ASAP7_75t_L g811 ( 
.A1(n_690),
.A2(n_600),
.A3(n_644),
.B(n_641),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_644),
.A2(n_641),
.B(n_634),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_645),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_720),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_666),
.B(n_539),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_644),
.A2(n_641),
.B(n_634),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_645),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_464),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_666),
.B(n_539),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_636),
.A2(n_561),
.B1(n_464),
.B2(n_676),
.Y(n_820)
);

AND3x2_ASAP7_75t_L g821 ( 
.A(n_704),
.B(n_575),
.C(n_362),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_539),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_730),
.B(n_731),
.Y(n_823)
);

AO21x1_ASAP7_75t_L g824 ( 
.A1(n_796),
.A2(n_737),
.B(n_805),
.Y(n_824)
);

NOR2x1_ASAP7_75t_SL g825 ( 
.A(n_778),
.B(n_780),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_795),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_781),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_793),
.B(n_785),
.Y(n_828)
);

BUFx2_ASAP7_75t_R g829 ( 
.A(n_798),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_815),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_819),
.B(n_822),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_766),
.A2(n_791),
.B(n_788),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_790),
.A2(n_812),
.B(n_807),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_808),
.Y(n_834)
);

OAI21x1_ASAP7_75t_SL g835 ( 
.A1(n_757),
.A2(n_741),
.B(n_736),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_784),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_816),
.A2(n_762),
.B(n_751),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_804),
.A2(n_820),
.B1(n_786),
.B2(n_738),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_743),
.B(n_800),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_782),
.B(n_789),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_742),
.A2(n_797),
.B(n_803),
.Y(n_841)
);

OAI21x1_ASAP7_75t_SL g842 ( 
.A1(n_777),
.A2(n_750),
.B(n_760),
.Y(n_842)
);

BUFx2_ASAP7_75t_SL g843 ( 
.A(n_748),
.Y(n_843)
);

AO222x2_ASAP7_75t_L g844 ( 
.A1(n_747),
.A2(n_749),
.B1(n_753),
.B2(n_818),
.C1(n_806),
.C2(n_801),
.Y(n_844)
);

AO21x2_ASAP7_75t_L g845 ( 
.A1(n_775),
.A2(n_746),
.B(n_734),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_779),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_814),
.B(n_754),
.Y(n_847)
);

AO31x2_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_758),
.A3(n_739),
.B(n_759),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_767),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_767),
.Y(n_850)
);

AO31x2_ASAP7_75t_L g851 ( 
.A1(n_792),
.A2(n_811),
.A3(n_809),
.B(n_745),
.Y(n_851)
);

OAI21x1_ASAP7_75t_SL g852 ( 
.A1(n_777),
.A2(n_769),
.B(n_771),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_802),
.A2(n_735),
.B(n_770),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_813),
.B(n_817),
.Y(n_854)
);

INVx11_ASAP7_75t_L g855 ( 
.A(n_767),
.Y(n_855)
);

CKINVDCx16_ASAP7_75t_R g856 ( 
.A(n_740),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_773),
.A2(n_768),
.B(n_764),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_792),
.A2(n_809),
.B(n_811),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_761),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_733),
.B(n_732),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_763),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_744),
.B(n_761),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_821),
.Y(n_863)
);

INVx4_ASAP7_75t_SL g864 ( 
.A(n_767),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_756),
.B(n_733),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_SL g866 ( 
.A1(n_787),
.A2(n_794),
.B(n_799),
.Y(n_866)
);

AO31x2_ASAP7_75t_L g867 ( 
.A1(n_745),
.A2(n_729),
.A3(n_776),
.B(n_756),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_755),
.A2(n_756),
.B(n_745),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_774),
.A2(n_729),
.B(n_776),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_729),
.A2(n_776),
.B(n_765),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_738),
.B(n_687),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_793),
.B(n_783),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_752),
.Y(n_873)
);

BUFx12f_ASAP7_75t_L g874 ( 
.A(n_747),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_795),
.Y(n_875)
);

AOI21xp33_ASAP7_75t_SL g876 ( 
.A1(n_795),
.A2(n_545),
.B(n_708),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_795),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_783),
.B(n_595),
.Y(n_878)
);

AO21x2_ASAP7_75t_L g879 ( 
.A1(n_790),
.A2(n_812),
.B(n_807),
.Y(n_879)
);

BUFx4f_ASAP7_75t_L g880 ( 
.A(n_738),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_730),
.Y(n_881)
);

NAND2x1p5_ASAP7_75t_L g882 ( 
.A(n_738),
.B(n_687),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_752),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_865),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_865),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_864),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_870),
.A2(n_841),
.B(n_832),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_878),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_825),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_830),
.B(n_831),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_842),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_850),
.B(n_827),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_879),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_879),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_864),
.B(n_849),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_837),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_873),
.B(n_883),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_864),
.B(n_853),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_880),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_873),
.B(n_883),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_855),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_880),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_877),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_836),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_881),
.Y(n_908)
);

INVxp33_ASAP7_75t_L g909 ( 
.A(n_840),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_871),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_860),
.B(n_857),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_838),
.B(n_854),
.Y(n_912)
);

AO21x2_ASAP7_75t_L g913 ( 
.A1(n_870),
.A2(n_841),
.B(n_869),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_877),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_844),
.B(n_876),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_884),
.B(n_851),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_884),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_906),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_885),
.B(n_824),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_893),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_913),
.B(n_851),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_899),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_898),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_913),
.B(n_858),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_913),
.B(n_867),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_915),
.A2(n_838),
.B1(n_882),
.B2(n_871),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_907),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_SL g928 ( 
.A1(n_910),
.A2(n_882),
.B1(n_835),
.B2(n_856),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_889),
.A2(n_863),
.B(n_828),
.C(n_872),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_902),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_901),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_900),
.B(n_867),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_892),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_901),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_894),
.B(n_868),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_900),
.B(n_868),
.Y(n_936)
);

NAND2x1_ASAP7_75t_L g937 ( 
.A(n_901),
.B(n_852),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_895),
.B(n_845),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_889),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_939),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_922),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_R g942 ( 
.A(n_939),
.B(n_902),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_927),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_922),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_916),
.B(n_921),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_916),
.B(n_887),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_923),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_927),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_931),
.B(n_934),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_920),
.B(n_886),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_916),
.B(n_921),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_936),
.B(n_903),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_921),
.B(n_887),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_933),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_917),
.B(n_903),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_918),
.B(n_844),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_925),
.B(n_935),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_936),
.B(n_890),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_925),
.B(n_887),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_933),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_931),
.B(n_911),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_945),
.B(n_924),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_945),
.B(n_924),
.Y(n_963)
);

NOR3x1_ASAP7_75t_L g964 ( 
.A(n_952),
.B(n_905),
.C(n_904),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_957),
.B(n_919),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_943),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_951),
.B(n_924),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_941),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_951),
.B(n_932),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_957),
.B(n_932),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_941),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_943),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_952),
.B(n_919),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_949),
.B(n_931),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_948),
.B(n_958),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_947),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_949),
.B(n_934),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_948),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_944),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_946),
.B(n_925),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_946),
.B(n_938),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_962),
.B(n_953),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_964),
.B(n_950),
.Y(n_983)
);

NAND4xp25_ASAP7_75t_L g984 ( 
.A(n_973),
.B(n_926),
.C(n_956),
.D(n_928),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_980),
.B(n_953),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_966),
.A2(n_910),
.B(n_920),
.C(n_909),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_962),
.B(n_959),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_969),
.B(n_958),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_975),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_972),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_976),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_980),
.B(n_959),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_974),
.A2(n_928),
.B(n_926),
.C(n_940),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_974),
.B(n_940),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_969),
.B(n_955),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_974),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_970),
.B(n_955),
.Y(n_997)
);

NAND4xp25_ASAP7_75t_L g998 ( 
.A(n_973),
.B(n_942),
.C(n_912),
.D(n_914),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_978),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_963),
.B(n_961),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_982),
.B(n_963),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_991),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_983),
.A2(n_970),
.B1(n_930),
.B2(n_950),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_991),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_988),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_989),
.B(n_967),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_995),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_983),
.A2(n_993),
.B1(n_994),
.B2(n_996),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_990),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_997),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_993),
.A2(n_905),
.B(n_920),
.C(n_950),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_998),
.B(n_829),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_985),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_SL g1015 ( 
.A1(n_984),
.A2(n_977),
.B(n_896),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_994),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_874),
.Y(n_1017)
);

OAI32xp33_ASAP7_75t_L g1018 ( 
.A1(n_1008),
.A2(n_930),
.A3(n_996),
.B1(n_940),
.B2(n_975),
.Y(n_1018)
);

OAI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_1013),
.A2(n_1015),
.B1(n_1003),
.B2(n_1016),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1014),
.B(n_982),
.Y(n_1020)
);

AOI222xp33_ASAP7_75t_L g1021 ( 
.A1(n_1012),
.A2(n_908),
.B1(n_897),
.B2(n_967),
.C1(n_987),
.C2(n_965),
.Y(n_1021)
);

OAI32xp33_ASAP7_75t_L g1022 ( 
.A1(n_1007),
.A2(n_1000),
.A3(n_910),
.B1(n_987),
.B2(n_954),
.Y(n_1022)
);

AOI322xp5_ASAP7_75t_L g1023 ( 
.A1(n_1005),
.A2(n_1000),
.A3(n_981),
.B1(n_977),
.B2(n_960),
.C1(n_954),
.C2(n_891),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1005),
.B(n_981),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1009),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_1018),
.A2(n_1012),
.B(n_1016),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_1019),
.A2(n_1017),
.B1(n_1010),
.B2(n_1011),
.C(n_1006),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_1022),
.A2(n_929),
.B(n_937),
.C(n_986),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_1021),
.A2(n_920),
.B(n_1002),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1025),
.B(n_1001),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_1020),
.A2(n_823),
.B(n_846),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_1024),
.A2(n_1004),
.B(n_1002),
.C(n_937),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1023),
.A2(n_1001),
.B1(n_1004),
.B2(n_888),
.C(n_979),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1033),
.B(n_968),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_1027),
.B(n_826),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1031),
.B(n_829),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_968),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_971),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1032),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_1035),
.B(n_843),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1034),
.B(n_1026),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_1036),
.B(n_875),
.C(n_826),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_1037),
.B(n_834),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_1039),
.B(n_1028),
.C(n_1038),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_SL g1045 ( 
.A(n_1039),
.B(n_875),
.C(n_840),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1040),
.B(n_834),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1043),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_1045),
.B(n_866),
.C(n_859),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1042),
.B(n_823),
.Y(n_1049)
);

NAND4xp75_ASAP7_75t_L g1050 ( 
.A(n_1041),
.B(n_904),
.C(n_862),
.D(n_823),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1047),
.B(n_1044),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_1049),
.B(n_859),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_L g1053 ( 
.A1(n_1051),
.A2(n_1046),
.B1(n_1052),
.B2(n_1050),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1053),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_1054),
.B(n_1048),
.C(n_847),
.Y(n_1055)
);

INVxp33_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1056),
.B(n_1050),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_1057),
.B(n_847),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_SL g1059 ( 
.A1(n_1058),
.A2(n_847),
.B1(n_861),
.B2(n_910),
.Y(n_1059)
);


endmodule