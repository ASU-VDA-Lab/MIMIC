module real_jpeg_32842_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_1),
.A2(n_213),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_1),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_1),
.A2(n_231),
.B1(n_261),
.B2(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_1),
.A2(n_231),
.B1(n_367),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_1),
.A2(n_231),
.B1(n_512),
.B2(n_514),
.Y(n_511)
);

OAI22x1_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_2),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_2),
.A2(n_147),
.B1(n_213),
.B2(n_218),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_2),
.A2(n_147),
.B1(n_441),
.B2(n_443),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_2),
.A2(n_147),
.B1(n_548),
.B2(n_553),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_4),
.A2(n_88),
.B1(n_232),
.B2(n_456),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_4),
.A2(n_88),
.B1(n_536),
.B2(n_540),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_5),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_5),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_5),
.A2(n_452),
.B1(n_529),
.B2(n_532),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_6),
.A2(n_121),
.B1(n_125),
.B2(n_130),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_130),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_6),
.A2(n_130),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_6),
.A2(n_130),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_7),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_7),
.A2(n_115),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_7),
.A2(n_115),
.B1(n_214),
.B2(n_353),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_7),
.A2(n_115),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_192),
.B1(n_193),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_8),
.A2(n_192),
.B1(n_241),
.B2(n_245),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_8),
.A2(n_192),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_8),
.A2(n_192),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_10),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_57),
.B(n_170),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_10),
.A2(n_137),
.A3(n_250),
.B1(n_253),
.B2(n_256),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_10),
.A2(n_64),
.B1(n_278),
.B2(n_284),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_10),
.B(n_349),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_10),
.A2(n_158),
.B1(n_366),
.B2(n_369),
.Y(n_365)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_13),
.Y(n_206)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_13),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_16),
.A2(n_424),
.B(n_426),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_16),
.B(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_16),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_16),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_17),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_17),
.A2(n_70),
.B1(n_414),
.B2(n_417),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_17),
.A2(n_70),
.B1(n_501),
.B2(n_504),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_18),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_18),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_19),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_19),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_517),
.Y(n_24)
);

OAI21x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_475),
.B(n_515),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_385),
.B(n_472),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_271),
.B(n_384),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_234),
.Y(n_29)
);

NOR2xp67_ASAP7_75t_SL g384 ( 
.A(n_30),
.B(n_234),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_167),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_94),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_32),
.B(n_94),
.C(n_167),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_62),
.B1(n_92),
.B2(n_93),
.Y(n_32)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_33),
.B(n_93),
.Y(n_396)
);

OAI32xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.A3(n_42),
.B1(n_48),
.B2(n_56),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_37),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_41),
.Y(n_180)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_45),
.Y(n_555)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_47),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_54),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_61),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_61),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_61),
.Y(n_514)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_79),
.B2(n_82),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_69),
.B1(n_143),
.B2(n_153),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_63),
.A2(n_143),
.B1(n_260),
.B2(n_269),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_63),
.A2(n_79),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_63),
.B(n_82),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_63),
.A2(n_79),
.B(n_449),
.Y(n_486)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_64),
.A2(n_278),
.B1(n_295),
.B2(n_302),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_64),
.A2(n_335),
.B1(n_344),
.B2(n_346),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_64),
.A2(n_423),
.B(n_448),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_66),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_66),
.Y(n_422)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_67),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_68),
.Y(n_264)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_68),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_75),
.Y(n_453)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_78),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_79),
.B(n_449),
.Y(n_448)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_87),
.Y(n_292)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_91),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_141),
.C(n_157),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_95),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_110),
.B1(n_120),
.B2(n_131),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_96),
.A2(n_110),
.B1(n_131),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_96),
.A2(n_131),
.B1(n_191),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_97),
.Y(n_372)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_98),
.Y(n_349)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_105),
.B2(n_108),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_104),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_104),
.Y(n_229)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_106),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g458 ( 
.A(n_107),
.Y(n_458)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_113),
.Y(n_395)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_120),
.A2(n_131),
.B1(n_365),
.B2(n_372),
.Y(n_364)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_123),
.Y(n_442)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_124),
.Y(n_541)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_129),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_131),
.A2(n_372),
.B1(n_392),
.B2(n_440),
.Y(n_439)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_137),
.B(n_140),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_132),
.A2(n_137),
.B(n_140),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_161),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_139),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_139),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_141),
.A2(n_142),
.B1(n_157),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_146),
.Y(n_301)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_152),
.Y(n_425)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_158),
.B(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_158),
.B(n_201),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_158),
.A2(n_253),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_158),
.B(n_318),
.Y(n_317)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_169),
.B1(n_172),
.B2(n_183),
.Y(n_168)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_159),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_159),
.A2(n_172),
.B1(n_402),
.B2(n_431),
.Y(n_430)
);

OAI22x1_ASAP7_75t_L g509 ( 
.A1(n_159),
.A2(n_172),
.B1(n_431),
.B2(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_159),
.B(n_559),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_163),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_166),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_189),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_168),
.B(n_190),
.C(n_200),
.Y(n_465)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_172),
.Y(n_399)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_173),
.B(n_511),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_177),
.Y(n_408)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_178),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_178),
.Y(n_434)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_178),
.Y(n_438)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_178),
.Y(n_552)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_183),
.Y(n_398)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_195),
.Y(n_444)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_212),
.B1(n_221),
.B2(n_230),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_221),
.B1(n_230),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_201),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_201),
.A2(n_221),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_201),
.A2(n_212),
.B1(n_221),
.B2(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_201),
.A2(n_221),
.B1(n_413),
.B2(n_455),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_201),
.A2(n_221),
.B1(n_455),
.B2(n_489),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_222),
.B(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_207),
.B1(n_209),
.B2(n_211),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_206),
.Y(n_327)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_220),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_221),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_222),
.Y(n_331)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_248),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_235),
.B(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_238),
.B(n_248),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_240),
.A2(n_315),
.B1(n_320),
.B2(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_241),
.Y(n_490)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_247),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_249),
.A2(n_258),
.B1(n_259),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_249),
.Y(n_362)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_260),
.Y(n_346)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_263),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx4f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_379),
.B(n_383),
.Y(n_271)
);

OAI31xp67_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_357),
.A3(n_377),
.B(n_378),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_339),
.B(n_340),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_305),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_293),
.B(n_304),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_303),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_301),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_332),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_332),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_321),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_R g341 ( 
.A(n_307),
.B(n_321),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_315),
.B1(n_316),
.B2(n_320),
.Y(n_307)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_310),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_315),
.A2(n_320),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AO22x1_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_328),
.B1(n_329),
.B2(n_331),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_342),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_355),
.C(n_359),
.Y(n_358)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_355),
.B2(n_356),
.Y(n_347)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_348),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_349),
.A2(n_500),
.B1(n_507),
.B2(n_508),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_349),
.A2(n_500),
.B1(n_508),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_360),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_373),
.C(n_376),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_373),
.B1(n_375),
.B2(n_376),
.Y(n_363)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_380),
.B(n_381),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_466),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_459),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_388),
.B(n_459),
.C(n_474),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_409),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_389),
.B(n_410),
.C(n_446),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_396),
.C(n_397),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_390),
.A2(n_391),
.B1(n_397),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

AOI22x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_400),
.A2(n_547),
.B(n_556),
.Y(n_546)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_445),
.Y(n_409)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_429),
.Y(n_410)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_420),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_420),
.Y(n_464)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_423),
.B(n_428),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_439),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g483 ( 
.A(n_439),
.Y(n_483)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_454),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.C(n_465),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_470),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_463),
.A2(n_464),
.B1(n_465),
.B2(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_465),
.Y(n_471)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_469),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_479),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_485),
.C(n_496),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_496),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_495),
.Y(n_485)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_486),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_486),
.B(n_488),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_489),
.Y(n_526)
);

BUFx6f_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_495),
.A2(n_546),
.B1(n_558),
.B2(n_560),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_495),
.B(n_557),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_509),
.C(n_522),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_509),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx4_ASAP7_75t_SL g512 ( 
.A(n_513),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_561),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_519),
.B(n_520),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_543),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_534),
.B(n_542),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_534),
.Y(n_542)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx3_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_547),
.Y(n_559)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);


endmodule