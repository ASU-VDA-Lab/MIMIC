module fake_jpeg_18959_n_33 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_23),
.B1(n_15),
.B2(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_22),
.B1(n_18),
.B2(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_5),
.Y(n_30)
);

AOI21x1_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_6),
.B(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_20),
.Y(n_33)
);


endmodule