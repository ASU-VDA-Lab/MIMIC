module fake_aes_7908_n_1374 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1374);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1374;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g301 ( .A(n_34), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_223), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_282), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_85), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_218), .Y(n_305) );
INVxp33_ASAP7_75t_L g306 ( .A(n_128), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_295), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_108), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_169), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_248), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_52), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_233), .Y(n_312) );
INVxp33_ASAP7_75t_SL g313 ( .A(n_274), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_0), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_13), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_289), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_88), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_249), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_220), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_148), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_104), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_36), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_38), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_47), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_73), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_266), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_96), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_141), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_152), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_151), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_176), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_103), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_77), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_149), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_213), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_1), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_203), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_48), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_48), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_262), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_45), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_263), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_30), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_278), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_25), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_66), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_280), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_71), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_250), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_30), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_102), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_26), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_2), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_62), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_75), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_90), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_118), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_114), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_276), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_243), .Y(n_362) );
BUFx10_ASAP7_75t_L g363 ( .A(n_26), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_54), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_230), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_36), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_86), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_166), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_83), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_60), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_159), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_154), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_42), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_76), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_14), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_290), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_21), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_300), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_299), .Y(n_379) );
BUFx10_ASAP7_75t_L g380 ( .A(n_127), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_283), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_49), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_109), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_78), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_94), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_15), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_201), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_116), .Y(n_388) );
INVxp33_ASAP7_75t_L g389 ( .A(n_56), .Y(n_389) );
INVxp33_ASAP7_75t_SL g390 ( .A(n_185), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_222), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_87), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_98), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_3), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_229), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_247), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_293), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_8), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_191), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_246), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_57), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_245), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_49), .Y(n_403) );
INVxp33_ASAP7_75t_SL g404 ( .A(n_133), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_63), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_135), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_13), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_129), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_22), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_270), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_93), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_193), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_180), .B(n_208), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_137), .Y(n_414) );
INVxp33_ASAP7_75t_SL g415 ( .A(n_158), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_297), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_111), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_165), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_195), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_164), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_61), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_63), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_237), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_175), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_147), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_288), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_107), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_38), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_255), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_35), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_272), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_285), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_162), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_186), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_173), .Y(n_435) );
INVxp33_ASAP7_75t_L g436 ( .A(n_50), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_3), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_51), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_194), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_252), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_296), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_46), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_235), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_95), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_142), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_273), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_8), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_19), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_227), .Y(n_449) );
INVx4_ASAP7_75t_L g450 ( .A(n_373), .Y(n_450) );
XOR2xp5_ASAP7_75t_L g451 ( .A(n_346), .B(n_0), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_389), .B(n_1), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_373), .Y(n_453) );
NAND2xp33_ASAP7_75t_L g454 ( .A(n_306), .B(n_69), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_402), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_317), .B(n_2), .Y(n_456) );
INVxp33_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_322), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_335), .Y(n_459) );
AND2x6_ASAP7_75t_L g460 ( .A(n_337), .B(n_70), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_335), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_303), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_322), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_303), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_353), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_380), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_436), .B(n_426), .Y(n_467) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_325), .A2(n_74), .B(n_72), .Y(n_468) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_325), .B(n_79), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_436), .B(n_4), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_335), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_301), .B(n_4), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_422), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_341), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_306), .B(n_5), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_341), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_347), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_380), .Y(n_478) );
CKINVDCx8_ASAP7_75t_R g479 ( .A(n_318), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_380), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_335), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_351), .Y(n_483) );
NOR2xp33_ASAP7_75t_SL g484 ( .A(n_318), .B(n_298), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_466), .B(n_347), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_460), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_475), .B(n_405), .C(n_351), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
INVx4_ASAP7_75t_SL g489 ( .A(n_460), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_453), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_473), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_466), .B(n_405), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_466), .B(n_333), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_483), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_466), .B(n_428), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_479), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_428), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_467), .B(n_438), .Y(n_500) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_457), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_478), .B(n_438), .Y(n_502) );
INVx5_ASAP7_75t_L g503 ( .A(n_460), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_457), .A2(n_315), .B1(n_307), .B2(n_305), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_469), .B(n_359), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_467), .A2(n_315), .B1(n_448), .B2(n_346), .Y(n_506) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_454), .A2(n_309), .B(n_302), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_450), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_452), .A2(n_311), .B1(n_324), .B2(n_323), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_470), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_478), .B(n_372), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_469), .B(n_359), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_470), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_470), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_465), .A2(n_448), .B1(n_403), .B2(n_305), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_459), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_478), .B(n_361), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_478), .Y(n_521) );
AO22x2_ASAP7_75t_L g522 ( .A1(n_456), .A2(n_355), .B1(n_338), .B2(n_339), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_451), .B(n_336), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
AND2x6_ASAP7_75t_L g527 ( .A(n_456), .B(n_337), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_469), .A2(n_364), .B1(n_366), .B2(n_354), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g529 ( .A(n_460), .B(n_423), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_456), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_491), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_495), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_522), .A2(n_469), .B1(n_456), .B2(n_454), .Y(n_534) );
OR2x6_ASAP7_75t_L g535 ( .A(n_504), .B(n_524), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_486), .B(n_479), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_493), .B(n_480), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_501), .B(n_480), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_499), .B(n_456), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_485), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_491), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_512), .B(n_465), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_485), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_522), .A2(n_475), .B1(n_484), .B2(n_472), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_522), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_500), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_492), .B(n_480), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_528), .A2(n_484), .B1(n_472), .B2(n_390), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_506), .B(n_464), .C(n_462), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_515), .B(n_307), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_496), .B(n_479), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_521), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_486), .B(n_455), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_498), .B(n_450), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_527), .Y(n_557) );
AND2x6_ASAP7_75t_L g558 ( .A(n_530), .B(n_383), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_486), .B(n_412), .Y(n_559) );
NOR3xp33_ASAP7_75t_SL g560 ( .A(n_517), .B(n_343), .C(n_314), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_488), .B(n_363), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_527), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_502), .B(n_450), .Y(n_563) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_520), .B(n_316), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_494), .B(n_450), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
OAI22xp5_ASAP7_75t_SL g567 ( .A1(n_525), .A2(n_451), .B1(n_473), .B2(n_316), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_494), .B(n_313), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_527), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_497), .A2(n_345), .B1(n_387), .B2(n_374), .Y(n_570) );
INVx5_ASAP7_75t_L g571 ( .A(n_527), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_527), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_520), .B(n_370), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_490), .B(n_313), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_519), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_511), .A2(n_374), .B1(n_387), .B2(n_345), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_513), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_505), .B(n_412), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_497), .B(n_416), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_487), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_503), .B(n_416), .Y(n_585) );
NAND2xp33_ASAP7_75t_SL g586 ( .A(n_505), .B(n_399), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_510), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_514), .A2(n_404), .B1(n_415), .B2(n_390), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_507), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_514), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_529), .A2(n_463), .B(n_474), .C(n_458), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_523), .B(n_420), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_489), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_503), .Y(n_595) );
INVx5_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_523), .B(n_404), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_489), .B(n_420), .Y(n_598) );
AND3x1_ASAP7_75t_L g599 ( .A(n_508), .B(n_377), .C(n_375), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_503), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_508), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_503), .B(n_432), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_489), .Y(n_603) );
AND2x6_ASAP7_75t_L g604 ( .A(n_529), .B(n_383), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_509), .B(n_447), .Y(n_605) );
AND2x6_ASAP7_75t_L g606 ( .A(n_509), .B(n_419), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_518), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_495), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_493), .B(n_399), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_495), .Y(n_611) );
AND2x6_ASAP7_75t_L g612 ( .A(n_530), .B(n_419), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_522), .A2(n_415), .B1(n_460), .B2(n_382), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_486), .B(n_432), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_500), .B(n_458), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_495), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_505), .A2(n_468), .B(n_368), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_555), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_596), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_596), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_609), .B(n_363), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_611), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_533), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_580), .B(n_443), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_578), .A2(n_443), .B1(n_386), .B2(n_398), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_546), .B(n_363), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_545), .A2(n_460), .B1(n_394), .B2(n_407), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_616), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_532), .Y(n_629) );
CKINVDCx11_ASAP7_75t_R g630 ( .A(n_535), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_557), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_571), .Y(n_632) );
INVx5_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
BUFx5_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_581), .B(n_401), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_566), .B(n_409), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_550), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_577), .B(n_421), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_541), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_537), .B(n_430), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_537), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_596), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_575), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_590), .B(n_437), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_540), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_531), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx4_ASAP7_75t_L g648 ( .A(n_571), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_573), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_592), .Y(n_650) );
INVx3_ASAP7_75t_L g651 ( .A(n_569), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_564), .B(n_433), .Y(n_652) );
AND2x4_ASAP7_75t_SL g653 ( .A(n_550), .B(n_610), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_534), .A2(n_442), .B(n_474), .C(n_463), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_543), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
CKINVDCx11_ASAP7_75t_R g657 ( .A(n_535), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_568), .B(n_355), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_578), .B(n_476), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_617), .A2(n_468), .B(n_312), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_607), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_542), .B(n_433), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_565), .A2(n_468), .B(n_332), .Y(n_663) );
OAI22x1_ASAP7_75t_L g664 ( .A1(n_610), .A2(n_365), .B1(n_304), .B2(n_468), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_553), .Y(n_665) );
BUFx10_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_607), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_615), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_568), .B(n_539), .Y(n_669) );
BUFx12f_ASAP7_75t_L g670 ( .A(n_535), .Y(n_670) );
BUFx12f_ASAP7_75t_L g671 ( .A(n_561), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_601), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_567), .B(n_476), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_570), .B(n_477), .Y(n_674) );
INVx3_ASAP7_75t_L g675 ( .A(n_569), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_605), .Y(n_676) );
BUFx8_ASAP7_75t_SL g677 ( .A(n_542), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_599), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_599), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_538), .B(n_477), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_539), .B(n_460), .Y(n_681) );
INVx3_ASAP7_75t_SL g682 ( .A(n_583), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_586), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_608), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_574), .A2(n_468), .B(n_368), .Y(n_685) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_564), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_589), .A2(n_319), .B(n_310), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_574), .Y(n_688) );
BUFx4f_ASAP7_75t_SL g689 ( .A(n_606), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_547), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_534), .A2(n_460), .B1(n_320), .B2(n_326), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_579), .Y(n_692) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_567), .A2(n_342), .B1(n_352), .B2(n_308), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_544), .A2(n_327), .B1(n_329), .B2(n_321), .Y(n_694) );
INVx4_ASAP7_75t_L g695 ( .A(n_558), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_613), .A2(n_460), .B1(n_330), .B2(n_334), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_556), .A2(n_340), .B(n_331), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_558), .Y(n_698) );
AND2x4_ASAP7_75t_SL g699 ( .A(n_549), .B(n_344), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_544), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_572), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_563), .A2(n_349), .B(n_348), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_548), .B(n_350), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_572), .B(n_369), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_595), .Y(n_705) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_572), .Y(n_706) );
BUFx3_ASAP7_75t_L g707 ( .A(n_606), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_554), .B(n_356), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_SL g709 ( .A1(n_576), .A2(n_413), .B(n_471), .C(n_461), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_548), .A2(n_357), .B1(n_360), .B2(n_358), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_588), .B(n_362), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_558), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_551), .B(n_367), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_560), .B(n_5), .Y(n_714) );
INVx1_ASAP7_75t_SL g715 ( .A(n_558), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_600), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_597), .B(n_6), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_L g718 ( .A1(n_591), .A2(n_378), .B(n_379), .C(n_376), .Y(n_718) );
BUFx12f_ASAP7_75t_L g719 ( .A(n_612), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_612), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_593), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_582), .B(n_328), .Y(n_722) );
INVxp67_ASAP7_75t_L g723 ( .A(n_612), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_598), .A2(n_384), .B1(n_393), .B2(n_388), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_612), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_606), .Y(n_726) );
NOR2xp33_ASAP7_75t_SL g727 ( .A(n_603), .B(n_396), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_606), .B(n_6), .Y(n_728) );
O2A1O1Ixp33_ASAP7_75t_L g729 ( .A1(n_559), .A2(n_391), .B(n_392), .C(n_381), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_594), .B(n_397), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_603), .B(n_439), .Y(n_731) );
OR2x6_ASAP7_75t_L g732 ( .A(n_536), .B(n_400), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_614), .Y(n_733) );
BUFx8_ASAP7_75t_L g734 ( .A(n_604), .Y(n_734) );
OR2x6_ASAP7_75t_L g735 ( .A(n_585), .B(n_406), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_602), .A2(n_445), .B1(n_446), .B2(n_440), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_604), .B(n_408), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_604), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_604), .Y(n_739) );
AOI21x1_ASAP7_75t_L g740 ( .A1(n_617), .A2(n_417), .B(n_410), .Y(n_740) );
CKINVDCx8_ASAP7_75t_R g741 ( .A(n_609), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_580), .A2(n_424), .B(n_425), .C(n_418), .Y(n_742) );
CKINVDCx11_ASAP7_75t_R g743 ( .A(n_532), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_609), .B(n_429), .Y(n_744) );
OAI21x1_ASAP7_75t_L g745 ( .A1(n_685), .A2(n_371), .B(n_361), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_618), .Y(n_746) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_741), .Y(n_747) );
AOI21x1_ASAP7_75t_L g748 ( .A1(n_740), .A2(n_385), .B(n_371), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_660), .A2(n_411), .B(n_385), .Y(n_749) );
OA21x2_ASAP7_75t_L g750 ( .A1(n_660), .A2(n_414), .B(n_411), .Y(n_750) );
AO21x2_ASAP7_75t_L g751 ( .A1(n_663), .A2(n_441), .B(n_431), .Y(n_751) );
NOR2xp67_ASAP7_75t_L g752 ( .A(n_623), .B(n_7), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_663), .A2(n_435), .B(n_414), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_672), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_668), .Y(n_755) );
OR2x2_ASAP7_75t_L g756 ( .A(n_622), .B(n_7), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_665), .Y(n_757) );
OR2x6_ASAP7_75t_L g758 ( .A(n_628), .B(n_435), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_669), .B(n_444), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_625), .A2(n_427), .B1(n_434), .B2(n_395), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_701), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_726), .A2(n_449), .B(n_461), .Y(n_762) );
OAI21x1_ASAP7_75t_L g763 ( .A1(n_738), .A2(n_471), .B(n_461), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g764 ( .A1(n_709), .A2(n_482), .B(n_481), .C(n_471), .Y(n_764) );
OR2x6_ASAP7_75t_L g765 ( .A(n_670), .B(n_427), .Y(n_765) );
INVx5_ASAP7_75t_L g766 ( .A(n_701), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_624), .B(n_9), .Y(n_767) );
BUFx2_ASAP7_75t_SL g768 ( .A(n_633), .Y(n_768) );
OAI21x1_ASAP7_75t_L g769 ( .A1(n_739), .A2(n_482), .B(n_481), .Y(n_769) );
OAI21x1_ASAP7_75t_L g770 ( .A1(n_725), .A2(n_482), .B(n_481), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_677), .Y(n_771) );
CKINVDCx6p67_ASAP7_75t_R g772 ( .A(n_743), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_687), .A2(n_423), .B(n_434), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_641), .Y(n_774) );
CKINVDCx16_ASAP7_75t_R g775 ( .A(n_671), .Y(n_775) );
AO21x2_ASAP7_75t_L g776 ( .A1(n_694), .A2(n_423), .B(n_81), .Y(n_776) );
AO31x2_ASAP7_75t_L g777 ( .A1(n_664), .A2(n_9), .A3(n_10), .B(n_11), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_640), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_629), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_669), .A2(n_10), .B(n_11), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_673), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_684), .Y(n_782) );
BUFx2_ASAP7_75t_R g783 ( .A(n_639), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_673), .A2(n_12), .B1(n_16), .B2(n_17), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_640), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_680), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_687), .A2(n_82), .B(n_80), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_624), .B(n_16), .Y(n_788) );
BUFx12f_ASAP7_75t_L g789 ( .A(n_630), .Y(n_789) );
AO31x2_ASAP7_75t_L g790 ( .A1(n_694), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_713), .A2(n_89), .B(n_84), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_648), .Y(n_792) );
OA21x2_ASAP7_75t_L g793 ( .A1(n_654), .A2(n_92), .B(n_91), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_702), .A2(n_18), .B(n_20), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_712), .A2(n_99), .B(n_97), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_656), .Y(n_796) );
OA21x2_ASAP7_75t_L g797 ( .A1(n_691), .A2(n_101), .B(n_100), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_690), .B(n_20), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_676), .B(n_21), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_712), .A2(n_106), .B(n_105), .Y(n_800) );
NOR2x1_ASAP7_75t_SL g801 ( .A(n_719), .B(n_22), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_688), .B(n_23), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_688), .B(n_23), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_692), .A2(n_112), .B(n_110), .Y(n_804) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_737), .A2(n_115), .B(n_113), .Y(n_805) );
AO31x2_ASAP7_75t_L g806 ( .A1(n_742), .A2(n_24), .A3(n_25), .B(n_27), .Y(n_806) );
AND2x4_ASAP7_75t_L g807 ( .A(n_695), .B(n_24), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_702), .A2(n_27), .B(n_28), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_700), .A2(n_28), .B1(n_29), .B2(n_31), .Y(n_809) );
AND2x4_ASAP7_75t_L g810 ( .A(n_695), .B(n_29), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_648), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_680), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g813 ( .A1(n_718), .A2(n_31), .B(n_32), .C(n_33), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_679), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_678), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_713), .A2(n_119), .B(n_117), .Y(n_816) );
OA21x2_ASAP7_75t_L g817 ( .A1(n_737), .A2(n_121), .B(n_120), .Y(n_817) );
OA21x2_ASAP7_75t_L g818 ( .A1(n_697), .A2(n_123), .B(n_122), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_710), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_653), .B(n_35), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_643), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_734), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_727), .B(n_37), .Y(n_823) );
AND2x4_ASAP7_75t_L g824 ( .A(n_646), .B(n_37), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_657), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_651), .A2(n_184), .B(n_292), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_621), .Y(n_827) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_661), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_734), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_655), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_647), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_645), .Y(n_832) );
INVx1_ASAP7_75t_SL g833 ( .A(n_701), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_SL g834 ( .A1(n_715), .A2(n_183), .B(n_291), .C(n_286), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_650), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_637), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_667), .Y(n_837) );
O2A1O1Ixp5_ASAP7_75t_L g838 ( .A1(n_686), .A2(n_182), .B(n_284), .C(n_281), .Y(n_838) );
OAI21x1_ASAP7_75t_L g839 ( .A1(n_651), .A2(n_179), .B(n_279), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_636), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_721), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_662), .B(n_39), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_658), .A2(n_178), .B(n_277), .Y(n_843) );
OAI21x1_ASAP7_75t_L g844 ( .A1(n_675), .A2(n_177), .B(n_275), .Y(n_844) );
OAI21x1_ASAP7_75t_L g845 ( .A1(n_675), .A2(n_642), .B(n_619), .Y(n_845) );
OAI22x1_ASAP7_75t_L g846 ( .A1(n_744), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_636), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_673), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_848) );
AO31x2_ASAP7_75t_L g849 ( .A1(n_703), .A2(n_43), .A3(n_44), .B(n_45), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_703), .A2(n_43), .B1(n_44), .B2(n_46), .Y(n_850) );
NOR2x1_ASAP7_75t_SL g851 ( .A(n_633), .B(n_47), .Y(n_851) );
AOI22x1_ASAP7_75t_L g852 ( .A1(n_717), .A2(n_681), .B1(n_697), .B2(n_733), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_635), .A2(n_638), .B1(n_658), .B2(n_693), .C(n_659), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_683), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_854) );
OR2x6_ASAP7_75t_L g855 ( .A(n_698), .B(n_53), .Y(n_855) );
A2O1A1Ixp33_ASAP7_75t_L g856 ( .A1(n_718), .A2(n_53), .B(n_54), .C(n_55), .Y(n_856) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_706), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_706), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_626), .B(n_682), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_619), .A2(n_196), .B(n_271), .Y(n_860) );
CKINVDCx14_ASAP7_75t_R g861 ( .A(n_714), .Y(n_861) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_706), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_644), .A2(n_192), .B(n_269), .Y(n_863) );
OAI21x1_ASAP7_75t_L g864 ( .A1(n_642), .A2(n_190), .B(n_268), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_638), .Y(n_865) );
OAI211xp5_ASAP7_75t_SL g866 ( .A1(n_674), .A2(n_55), .B(n_56), .C(n_57), .Y(n_866) );
INVxp67_ASAP7_75t_L g867 ( .A(n_728), .Y(n_867) );
AO21x2_ASAP7_75t_L g868 ( .A1(n_644), .A2(n_198), .B(n_267), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g869 ( .A(n_727), .B(n_58), .Y(n_869) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_627), .A2(n_197), .B(n_265), .Y(n_870) );
OAI21x1_ASAP7_75t_L g871 ( .A1(n_729), .A2(n_189), .B(n_264), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_666), .Y(n_872) );
AO31x2_ASAP7_75t_L g873 ( .A1(n_635), .A2(n_58), .A3(n_59), .B(n_60), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_696), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_874) );
A2O1A1Ixp33_ASAP7_75t_L g875 ( .A1(n_729), .A2(n_64), .B(n_65), .C(n_66), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_666), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_711), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_620), .A2(n_202), .B(n_261), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_681), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_633), .B(n_64), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g881 ( .A(n_633), .B(n_65), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_715), .A2(n_67), .B1(n_68), .B2(n_124), .Y(n_882) );
O2A1O1Ixp33_ASAP7_75t_L g883 ( .A1(n_711), .A2(n_67), .B(n_68), .C(n_125), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_853), .A2(n_699), .B1(n_722), .B2(n_708), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_761), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_840), .A2(n_847), .B1(n_865), .B2(n_848), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_841), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_853), .B(n_730), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_767), .A2(n_708), .B1(n_730), .B2(n_652), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_877), .B(n_732), .Y(n_890) );
INVx5_ASAP7_75t_SL g891 ( .A(n_772), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_827), .A2(n_732), .B1(n_735), .B2(n_689), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_775), .B(n_705), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_842), .A2(n_732), .B1(n_735), .B2(n_704), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_824), .A2(n_735), .B1(n_716), .B2(n_707), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_766), .Y(n_896) );
AOI222xp33_ASAP7_75t_L g897 ( .A1(n_755), .A2(n_723), .B1(n_720), .B2(n_731), .C1(n_724), .C2(n_632), .Y(n_897) );
NAND2xp5_ASAP7_75t_SL g898 ( .A(n_807), .B(n_631), .Y(n_898) );
CKINVDCx6p67_ASAP7_75t_R g899 ( .A(n_747), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_824), .A2(n_632), .B1(n_634), .B2(n_649), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_753), .A2(n_649), .B(n_736), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_754), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_848), .A2(n_631), .B1(n_634), .B2(n_131), .Y(n_903) );
OAI21xp33_ASAP7_75t_SL g904 ( .A1(n_855), .A2(n_634), .B(n_631), .Y(n_904) );
INVxp67_ASAP7_75t_L g905 ( .A(n_802), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_746), .B(n_634), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_782), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_872), .B(n_876), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_757), .Y(n_909) );
O2A1O1Ixp33_ASAP7_75t_L g910 ( .A1(n_866), .A2(n_634), .B(n_130), .C(n_132), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_867), .A2(n_126), .B1(n_134), .B2(n_136), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_802), .B(n_138), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_758), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_756), .B(n_139), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_749), .A2(n_140), .B(n_143), .Y(n_915) );
AOI21x1_ASAP7_75t_L g916 ( .A1(n_748), .A2(n_144), .B(n_145), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_867), .A2(n_146), .B1(n_150), .B2(n_153), .Y(n_917) );
INVx5_ASAP7_75t_L g918 ( .A(n_761), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_796), .Y(n_919) );
BUFx3_ASAP7_75t_L g920 ( .A(n_771), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_830), .Y(n_921) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_761), .Y(n_922) );
AOI21x1_ASAP7_75t_L g923 ( .A1(n_750), .A2(n_155), .B(n_156), .Y(n_923) );
OAI211xp5_ASAP7_75t_L g924 ( .A1(n_819), .A2(n_157), .B(n_160), .C(n_161), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_798), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_778), .A2(n_163), .B1(n_167), .B2(n_168), .C(n_170), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_798), .Y(n_927) );
BUFx8_ASAP7_75t_SL g928 ( .A(n_789), .Y(n_928) );
BUFx2_ASAP7_75t_L g929 ( .A(n_758), .Y(n_929) );
AND2x6_ASAP7_75t_L g930 ( .A(n_807), .B(n_171), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_786), .B(n_294), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_759), .B(n_172), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_832), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_774), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_859), .A2(n_174), .B1(n_181), .B2(n_187), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_803), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_861), .A2(n_188), .B1(n_199), .B2(n_200), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_758), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_803), .Y(n_939) );
OA21x2_ASAP7_75t_L g940 ( .A1(n_745), .A2(n_204), .B(n_205), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_814), .B(n_206), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_855), .A2(n_207), .B1(n_209), .B2(n_210), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_850), .Y(n_943) );
NAND2x1_ASAP7_75t_L g944 ( .A(n_862), .B(n_211), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_759), .B(n_212), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_815), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_760), .A2(n_820), .B1(n_812), .B2(n_785), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_850), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_821), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_799), .A2(n_217), .B1(n_219), .B2(n_221), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_764), .A2(n_224), .B(n_225), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_788), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_879), .B(n_226), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_753), .A2(n_228), .B(n_231), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_855), .A2(n_232), .B1(n_234), .B2(n_236), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_809), .A2(n_238), .B1(n_239), .B2(n_240), .C(n_241), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_819), .A2(n_242), .B1(n_244), .B2(n_251), .Y(n_957) );
OAI21xp5_ASAP7_75t_L g958 ( .A1(n_773), .A2(n_253), .B(n_254), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_809), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_765), .A2(n_256), .B1(n_257), .B2(n_258), .C(n_259), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_873), .Y(n_961) );
AND2x4_ASAP7_75t_L g962 ( .A(n_822), .B(n_829), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_750), .A2(n_751), .B(n_816), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_783), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_836), .A2(n_810), .B1(n_852), .B2(n_765), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_873), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_810), .A2(n_765), .B1(n_866), .B2(n_752), .Y(n_967) );
A2O1A1Ixp33_ASAP7_75t_L g968 ( .A1(n_780), .A2(n_794), .B(n_808), .C(n_883), .Y(n_968) );
OAI21xp5_ASAP7_75t_L g969 ( .A1(n_794), .A2(n_808), .B(n_780), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_873), .Y(n_970) );
OAI221xp5_ASAP7_75t_L g971 ( .A1(n_781), .A2(n_784), .B1(n_813), .B2(n_856), .C(n_875), .Y(n_971) );
AOI21xp33_ASAP7_75t_L g972 ( .A1(n_883), .A2(n_751), .B(n_776), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_801), .A2(n_851), .B1(n_880), .B2(n_874), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_874), .A2(n_880), .B1(n_846), .B2(n_828), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_828), .A2(n_837), .B1(n_779), .B2(n_869), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_825), .A2(n_882), .B1(n_823), .B2(n_837), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_831), .B(n_835), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_882), .A2(n_854), .B1(n_797), .B2(n_766), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_768), .B(n_790), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_881), .A2(n_863), .B1(n_791), .B2(n_843), .C(n_792), .Y(n_980) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_863), .A2(n_791), .B1(n_843), .B2(n_811), .C(n_792), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_777), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_811), .A2(n_776), .B1(n_797), .B2(n_793), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_793), .A2(n_766), .B1(n_870), .B2(n_857), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_783), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_790), .B(n_806), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_790), .B(n_806), .Y(n_987) );
AO22x1_ASAP7_75t_L g988 ( .A1(n_766), .A2(n_857), .B1(n_862), .B2(n_833), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_833), .Y(n_989) );
BUFx6f_ASAP7_75t_L g990 ( .A(n_862), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_806), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_818), .A2(n_870), .B1(n_817), .B2(n_858), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_849), .B(n_777), .Y(n_993) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_849), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_849), .B(n_777), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_845), .B(n_871), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_834), .A2(n_838), .B1(n_868), .B2(n_787), .C(n_805), .Y(n_997) );
AO21x2_ASAP7_75t_L g998 ( .A1(n_868), .A2(n_804), .B(n_762), .Y(n_998) );
INVx4_ASAP7_75t_L g999 ( .A(n_860), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_864), .B(n_826), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_839), .B(n_844), .Y(n_1001) );
OAI21x1_ASAP7_75t_L g1002 ( .A1(n_763), .A2(n_769), .B(n_770), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_795), .Y(n_1003) );
AOI21xp5_ASAP7_75t_L g1004 ( .A1(n_838), .A2(n_878), .B(n_800), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_840), .B(n_546), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_853), .A2(n_741), .B1(n_611), .B2(n_616), .C(n_609), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_755), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_841), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_755), .Y(n_1009) );
OAI21x1_ASAP7_75t_L g1010 ( .A1(n_745), .A2(n_749), .B(n_763), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1005), .B(n_959), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_918), .B(n_979), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_982), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_991), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_918), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_961), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_888), .B(n_884), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_966), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_913), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_915), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_923), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_902), .B(n_907), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_887), .B(n_1008), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_918), .B(n_885), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_918), .B(n_885), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_919), .B(n_949), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_970), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_943), .B(n_948), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_925), .B(n_927), .Y(n_1029) );
INVxp67_ASAP7_75t_SL g1030 ( .A(n_905), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_886), .A2(n_974), .B1(n_973), .B2(n_895), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1003), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_987), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1034 ( .A(n_886), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_921), .B(n_909), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_896), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_999), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_986), .B(n_933), .Y(n_1038) );
OA21x2_ASAP7_75t_L g1039 ( .A1(n_972), .A2(n_963), .B(n_1004), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_930), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_993), .Y(n_1041) );
AOI222xp33_ASAP7_75t_L g1042 ( .A1(n_1006), .A2(n_952), .B1(n_891), .B2(n_969), .C1(n_929), .C2(n_938), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_977), .B(n_1007), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_989), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_999), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_890), .Y(n_1046) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_930), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_995), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1009), .B(n_934), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_885), .B(n_922), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_906), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_947), .B(n_890), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_906), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_969), .B(n_896), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_912), .B(n_936), .Y(n_1055) );
OR2x6_ASAP7_75t_L g1056 ( .A(n_903), .B(n_988), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_940), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_994), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_939), .B(n_968), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_967), .B(n_898), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_976), .A2(n_971), .B1(n_889), .B2(n_894), .C(n_965), .Y(n_1061) );
HB1xp67_ASAP7_75t_L g1062 ( .A(n_908), .Y(n_1062) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_922), .B(n_990), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1001), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_914), .B(n_941), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_892), .B(n_893), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_975), .B(n_945), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_953), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_930), .B(n_945), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_940), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_908), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_930), .B(n_932), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_932), .B(n_942), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_903), .B(n_978), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_942), .B(n_955), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_953), .Y(n_1076) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_955), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_920), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_996), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_998), .Y(n_1080) );
A2O1A1Ixp33_ASAP7_75t_L g1081 ( .A1(n_910), .A2(n_956), .B(n_904), .C(n_924), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_922), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_990), .B(n_1000), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_900), .B(n_990), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_954), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_897), .B(n_962), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_954), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_901), .B(n_931), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_981), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_998), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_901), .B(n_897), .Y(n_1091) );
NOR2x1_ASAP7_75t_SL g1092 ( .A(n_978), .B(n_992), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_972), .B(n_983), .Y(n_1093) );
BUFx3_ASAP7_75t_L g1094 ( .A(n_962), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_891), .Y(n_1095) );
OA21x2_ASAP7_75t_L g1096 ( .A1(n_997), .A2(n_984), .B(n_992), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_980), .B(n_957), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_958), .B(n_1010), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_958), .B(n_937), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_1002), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_911), .B(n_917), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_935), .B(n_950), .Y(n_1102) );
NOR3xp33_ASAP7_75t_SL g1103 ( .A(n_964), .B(n_985), .C(n_960), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_916), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_946), .B(n_926), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_944), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_891), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_899), .B(n_951), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_928), .B(n_902), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_913), .Y(n_1110) );
INVx3_ASAP7_75t_L g1111 ( .A(n_885), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_991), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_991), .Y(n_1113) );
OAI211xp5_ASAP7_75t_L g1114 ( .A1(n_1042), .A2(n_1086), .B(n_1061), .C(n_1108), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_1038), .B(n_1041), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1032), .Y(n_1116) );
OAI221xp5_ASAP7_75t_L g1117 ( .A1(n_1031), .A2(n_1066), .B1(n_1011), .B2(n_1067), .C(n_1052), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1038), .B(n_1041), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1043), .B(n_1029), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1014), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1014), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1048), .B(n_1054), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_1091), .A2(n_1075), .B1(n_1017), .B2(n_1077), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1048), .B(n_1054), .Y(n_1124) );
AND3x1_ASAP7_75t_L g1125 ( .A(n_1103), .B(n_1091), .C(n_1075), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1112), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1059), .B(n_1028), .Y(n_1127) );
OAI31xp33_ASAP7_75t_L g1128 ( .A1(n_1060), .A2(n_1040), .A3(n_1047), .B(n_1067), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1059), .B(n_1028), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1033), .B(n_1049), .Y(n_1130) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_1058), .A2(n_1089), .A3(n_1065), .B1(n_1033), .B2(n_1027), .B3(n_1018), .Y(n_1131) );
NAND3xp33_ASAP7_75t_L g1132 ( .A(n_1058), .B(n_1044), .C(n_1060), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1112), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_1083), .B(n_1012), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1049), .B(n_1064), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1064), .B(n_1034), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1113), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1043), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1035), .B(n_1051), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1035), .B(n_1051), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_1046), .B(n_1053), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1073), .A2(n_1102), .B1(n_1105), .B2(n_1040), .Y(n_1142) );
OAI33xp33_ASAP7_75t_L g1143 ( .A1(n_1089), .A2(n_1065), .A3(n_1027), .B1(n_1018), .B2(n_1016), .B3(n_1113), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1029), .B(n_1022), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1053), .B(n_1016), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1022), .B(n_1026), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1074), .B(n_1012), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1013), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1090), .Y(n_1149) );
OR2x6_ASAP7_75t_L g1150 ( .A(n_1047), .B(n_1056), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1023), .B(n_1026), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1023), .B(n_1012), .Y(n_1152) );
OR2x6_ASAP7_75t_L g1153 ( .A(n_1056), .B(n_1074), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1012), .B(n_1083), .Y(n_1154) );
INVx3_ASAP7_75t_L g1155 ( .A(n_1050), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1083), .B(n_1092), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1083), .B(n_1092), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1088), .B(n_1073), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1019), .B(n_1110), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1088), .B(n_1069), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1069), .B(n_1072), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1055), .B(n_1078), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1055), .B(n_1030), .Y(n_1163) );
OAI321xp33_ASAP7_75t_L g1164 ( .A1(n_1056), .A2(n_1097), .A3(n_1093), .B1(n_1099), .B2(n_1102), .C(n_1085), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1072), .B(n_1090), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1068), .B(n_1076), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1093), .B(n_1071), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1062), .B(n_1094), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1079), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1094), .B(n_1036), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1068), .B(n_1076), .Y(n_1171) );
A2O1A1Ixp33_ASAP7_75t_SL g1172 ( .A1(n_1106), .A2(n_1111), .B(n_1045), .C(n_1037), .Y(n_1172) );
AND2x4_ASAP7_75t_L g1173 ( .A(n_1037), .B(n_1045), .Y(n_1173) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1050), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1082), .B(n_1080), .Y(n_1175) );
INVx4_ASAP7_75t_L g1176 ( .A(n_1024), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_1056), .Y(n_1177) );
OAI221xp5_ASAP7_75t_SL g1178 ( .A1(n_1097), .A2(n_1056), .B1(n_1099), .B2(n_1081), .C(n_1094), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1179 ( .A(n_1109), .B(n_1095), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1180 ( .A(n_1087), .B(n_1045), .C(n_1107), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1100), .Y(n_1181) );
NAND2xp5_ASAP7_75t_SL g1182 ( .A(n_1015), .B(n_1036), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1036), .B(n_1015), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1084), .B(n_1096), .Y(n_1184) );
OR2x6_ASAP7_75t_L g1185 ( .A(n_1098), .B(n_1084), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1096), .B(n_1063), .Y(n_1186) );
INVx3_ASAP7_75t_L g1187 ( .A(n_1173), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1138), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1116), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1130), .Y(n_1190) );
OAI322xp33_ASAP7_75t_L g1191 ( .A1(n_1117), .A2(n_1109), .A3(n_1106), .B1(n_1105), .B2(n_1101), .C1(n_1020), .C2(n_1070), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1130), .Y(n_1192) );
BUFx2_ASAP7_75t_L g1193 ( .A(n_1176), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1115), .B(n_1111), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1115), .B(n_1111), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1142), .A2(n_1101), .B1(n_1098), .B2(n_1096), .Y(n_1196) );
NAND2xp33_ASAP7_75t_SL g1197 ( .A(n_1177), .B(n_1098), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1160), .B(n_1039), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1122), .B(n_1039), .Y(n_1199) );
OAI21xp5_ASAP7_75t_L g1200 ( .A1(n_1114), .A2(n_1024), .B(n_1025), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1122), .B(n_1039), .Y(n_1201) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_1132), .B(n_1111), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1135), .B(n_1024), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1119), .B(n_1024), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1205 ( .A(n_1156), .B(n_1098), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1124), .B(n_1039), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1135), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1120), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1118), .B(n_1025), .Y(n_1209) );
AOI211xp5_ASAP7_75t_SL g1210 ( .A1(n_1178), .A2(n_1025), .B(n_1050), .C(n_1063), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1146), .B(n_1025), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1120), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1118), .B(n_1050), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1146), .B(n_1063), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1124), .B(n_1100), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_1156), .B(n_1063), .Y(n_1216) );
NAND2x1p5_ASAP7_75t_L g1217 ( .A(n_1183), .B(n_1057), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1158), .B(n_1057), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1139), .B(n_1021), .Y(n_1219) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_1172), .A2(n_1104), .B(n_1021), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1163), .B(n_1159), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1139), .B(n_1104), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1158), .B(n_1104), .Y(n_1223) );
NOR2xp33_ASAP7_75t_SL g1224 ( .A(n_1176), .B(n_1183), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1140), .B(n_1144), .Y(n_1225) );
INVx1_ASAP7_75t_SL g1226 ( .A(n_1162), .Y(n_1226) );
NAND2xp5_ASAP7_75t_SL g1227 ( .A(n_1164), .B(n_1125), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_1125), .A2(n_1123), .B1(n_1153), .B2(n_1150), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1140), .B(n_1129), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1127), .B(n_1129), .Y(n_1230) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_1134), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1121), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1152), .B(n_1151), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1127), .B(n_1161), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1161), .B(n_1165), .Y(n_1235) );
NAND2x1_ASAP7_75t_L g1236 ( .A(n_1150), .B(n_1153), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1166), .B(n_1171), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1166), .B(n_1171), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1165), .B(n_1184), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1152), .B(n_1136), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1184), .B(n_1154), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1121), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1154), .B(n_1175), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1176), .B(n_1134), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1134), .B(n_1159), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1126), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1126), .Y(n_1247) );
AND2x2_ASAP7_75t_SL g1248 ( .A(n_1177), .B(n_1134), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1136), .B(n_1133), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1133), .B(n_1137), .Y(n_1250) );
OR2x6_ASAP7_75t_L g1251 ( .A(n_1150), .B(n_1153), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1226), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1239), .B(n_1186), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1239), .B(n_1186), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1190), .B(n_1149), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1241), .B(n_1185), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1241), .B(n_1185), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1235), .B(n_1185), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1208), .Y(n_1259) );
INVx2_ASAP7_75t_SL g1260 ( .A(n_1193), .Y(n_1260) );
AND2x4_ASAP7_75t_L g1261 ( .A(n_1205), .B(n_1157), .Y(n_1261) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1189), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1192), .B(n_1149), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1235), .B(n_1185), .Y(n_1264) );
AND3x2_ASAP7_75t_L g1265 ( .A(n_1224), .B(n_1128), .C(n_1157), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1207), .B(n_1137), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1212), .Y(n_1267) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1189), .Y(n_1268) );
NAND2xp5_ASAP7_75t_SL g1269 ( .A(n_1227), .B(n_1180), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1221), .B(n_1179), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1199), .B(n_1167), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1198), .B(n_1185), .Y(n_1272) );
OAI21xp33_ASAP7_75t_L g1273 ( .A1(n_1227), .A2(n_1153), .B(n_1150), .Y(n_1273) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1199), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1198), .B(n_1153), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1232), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1201), .B(n_1206), .Y(n_1277) );
NAND4xp25_ASAP7_75t_L g1278 ( .A(n_1196), .B(n_1167), .C(n_1168), .D(n_1141), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1201), .B(n_1145), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1234), .B(n_1147), .Y(n_1280) );
A2O1A1Ixp33_ASAP7_75t_L g1281 ( .A1(n_1210), .A2(n_1182), .B(n_1141), .C(n_1168), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1234), .B(n_1147), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1242), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1206), .B(n_1145), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1249), .B(n_1169), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1188), .B(n_1169), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1223), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1243), .B(n_1175), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1229), .B(n_1150), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1243), .B(n_1173), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1246), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1230), .B(n_1148), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1218), .B(n_1215), .Y(n_1293) );
OAI221xp5_ASAP7_75t_SL g1294 ( .A1(n_1273), .A2(n_1196), .B1(n_1251), .B2(n_1233), .C(n_1240), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1280), .B(n_1221), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1274), .Y(n_1296) );
NAND3xp33_ASAP7_75t_L g1297 ( .A(n_1269), .B(n_1202), .C(n_1228), .Y(n_1297) );
AOI211xp5_ASAP7_75t_SL g1298 ( .A1(n_1273), .A2(n_1191), .B(n_1202), .C(n_1216), .Y(n_1298) );
O2A1O1Ixp5_ASAP7_75t_L g1299 ( .A1(n_1281), .A2(n_1236), .B(n_1131), .C(n_1197), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g1300 ( .A(n_1252), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1301 ( .A(n_1260), .Y(n_1301) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_1278), .A2(n_1200), .B1(n_1197), .B2(n_1231), .C(n_1251), .Y(n_1302) );
OAI21xp33_ASAP7_75t_L g1303 ( .A1(n_1278), .A2(n_1245), .B(n_1251), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1274), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1292), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_1270), .A2(n_1248), .B1(n_1251), .B2(n_1231), .Y(n_1306) );
OAI32xp33_ASAP7_75t_L g1307 ( .A1(n_1289), .A2(n_1209), .A3(n_1225), .B1(n_1204), .B2(n_1237), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1274), .B(n_1218), .Y(n_1308) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1262), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1259), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_1275), .A2(n_1248), .B1(n_1214), .B2(n_1203), .Y(n_1311) );
OAI221xp5_ASAP7_75t_SL g1312 ( .A1(n_1289), .A2(n_1213), .B1(n_1238), .B2(n_1194), .C(n_1195), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1253), .B(n_1215), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1262), .Y(n_1314) );
NAND3x2_ASAP7_75t_L g1315 ( .A(n_1261), .B(n_1244), .C(n_1205), .Y(n_1315) );
O2A1O1Ixp33_ASAP7_75t_L g1316 ( .A1(n_1260), .A2(n_1143), .B(n_1170), .C(n_1250), .Y(n_1316) );
NOR2x1_ASAP7_75t_L g1317 ( .A(n_1261), .B(n_1173), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_1275), .A2(n_1205), .B1(n_1211), .B2(n_1216), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1259), .Y(n_1319) );
NAND3xp33_ASAP7_75t_L g1320 ( .A(n_1265), .B(n_1219), .C(n_1222), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1267), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_1298), .A2(n_1279), .B1(n_1284), .B2(n_1271), .Y(n_1322) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1309), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1315), .A2(n_1320), .B1(n_1294), .B2(n_1318), .Y(n_1324) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_1316), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1310), .Y(n_1326) );
XNOR2x1_ASAP7_75t_L g1327 ( .A(n_1315), .B(n_1265), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1310), .Y(n_1328) );
INVxp67_ASAP7_75t_SL g1329 ( .A(n_1300), .Y(n_1329) );
AOI21xp33_ASAP7_75t_L g1330 ( .A1(n_1297), .A2(n_1286), .B(n_1263), .Y(n_1330) );
INVx2_ASAP7_75t_L g1331 ( .A(n_1309), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1319), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1305), .B(n_1277), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1313), .B(n_1282), .Y(n_1334) );
XOR2x2_ASAP7_75t_L g1335 ( .A(n_1295), .B(n_1264), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1319), .Y(n_1336) );
AOI21xp5_ASAP7_75t_L g1337 ( .A1(n_1299), .A2(n_1261), .B(n_1285), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1321), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1313), .B(n_1282), .Y(n_1339) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_1317), .B(n_1261), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1341 ( .A1(n_1322), .A2(n_1307), .B1(n_1303), .B2(n_1312), .C(n_1302), .Y(n_1341) );
NOR2x1_ASAP7_75t_L g1342 ( .A(n_1327), .B(n_1321), .Y(n_1342) );
OAI21xp5_ASAP7_75t_L g1343 ( .A1(n_1322), .A2(n_1301), .B(n_1307), .Y(n_1343) );
OAI221xp5_ASAP7_75t_L g1344 ( .A1(n_1324), .A2(n_1306), .B1(n_1311), .B2(n_1304), .C(n_1296), .Y(n_1344) );
OAI221xp5_ASAP7_75t_L g1345 ( .A1(n_1325), .A2(n_1304), .B1(n_1296), .B2(n_1271), .C(n_1277), .Y(n_1345) );
OAI21xp5_ASAP7_75t_L g1346 ( .A1(n_1337), .A2(n_1258), .B(n_1257), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_1330), .A2(n_1216), .B1(n_1272), .B2(n_1187), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1329), .B(n_1253), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1329), .A2(n_1279), .B(n_1284), .Y(n_1349) );
OAI32xp33_ASAP7_75t_L g1350 ( .A1(n_1334), .A2(n_1257), .A3(n_1256), .B1(n_1308), .B2(n_1287), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1326), .Y(n_1351) );
OAI211xp5_ASAP7_75t_L g1352 ( .A1(n_1342), .A2(n_1339), .B(n_1256), .C(n_1333), .Y(n_1352) );
AOI22xp5_ASAP7_75t_L g1353 ( .A1(n_1341), .A2(n_1340), .B1(n_1335), .B2(n_1336), .Y(n_1353) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_1344), .A2(n_1340), .B1(n_1338), .B2(n_1332), .Y(n_1354) );
AOI222xp33_ASAP7_75t_L g1355 ( .A1(n_1343), .A2(n_1328), .B1(n_1254), .B2(n_1266), .C1(n_1263), .C2(n_1255), .Y(n_1355) );
A2O1A1Ixp33_ASAP7_75t_L g1356 ( .A1(n_1346), .A2(n_1308), .B(n_1290), .C(n_1254), .Y(n_1356) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_1347), .A2(n_1290), .B1(n_1293), .B2(n_1287), .Y(n_1357) );
AOI21xp33_ASAP7_75t_SL g1358 ( .A1(n_1345), .A2(n_1331), .B(n_1323), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g1359 ( .A1(n_1352), .A2(n_1349), .B(n_1350), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1353), .B(n_1347), .Y(n_1360) );
NAND3xp33_ASAP7_75t_L g1361 ( .A(n_1355), .B(n_1351), .C(n_1348), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1357), .B(n_1287), .Y(n_1362) );
NOR3xp33_ASAP7_75t_L g1363 ( .A(n_1360), .B(n_1358), .C(n_1354), .Y(n_1363) );
XOR2xp5_ASAP7_75t_L g1364 ( .A(n_1361), .B(n_1359), .Y(n_1364) );
AOI221xp5_ASAP7_75t_L g1365 ( .A1(n_1362), .A2(n_1356), .B1(n_1267), .B2(n_1276), .C(n_1283), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1364), .B(n_1288), .Y(n_1366) );
INVx1_ASAP7_75t_SL g1367 ( .A(n_1363), .Y(n_1367) );
OAI22xp5_ASAP7_75t_SL g1368 ( .A1(n_1367), .A2(n_1365), .B1(n_1217), .B2(n_1291), .Y(n_1368) );
AOI22xp5_ASAP7_75t_L g1369 ( .A1(n_1366), .A2(n_1276), .B1(n_1291), .B2(n_1174), .Y(n_1369) );
AOI22xp5_ASAP7_75t_L g1370 ( .A1(n_1368), .A2(n_1155), .B1(n_1174), .B2(n_1314), .Y(n_1370) );
OAI222xp33_ASAP7_75t_L g1371 ( .A1(n_1369), .A2(n_1285), .B1(n_1217), .B2(n_1220), .C1(n_1247), .C2(n_1174), .Y(n_1371) );
AO221x1_ASAP7_75t_L g1372 ( .A1(n_1371), .A2(n_1155), .B1(n_1187), .B2(n_1268), .C(n_1181), .Y(n_1372) );
NAND2xp5_ASAP7_75t_SL g1373 ( .A(n_1372), .B(n_1370), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g1374 ( .A1(n_1373), .A2(n_1268), .B(n_1155), .Y(n_1374) );
endmodule