module real_jpeg_24828_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_178;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

INVx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_62),
.B1(n_83),
.B2(n_108),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_62),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_11),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_82),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_82),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_82),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_13),
.A2(n_69),
.B1(n_109),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_13),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_132),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_132),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_67),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_67),
.Y(n_238)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_15),
.B(n_76),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_40),
.C(n_54),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_15),
.B(n_151),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_156),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_15),
.B(n_28),
.C(n_45),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_15),
.A2(n_30),
.B(n_239),
.Y(n_269)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_16),
.Y(n_163)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_20),
.B(n_113),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_112),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.C(n_64),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_23),
.A2(n_24),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_25),
.A2(n_35),
.B1(n_36),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_25),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_26),
.A2(n_30),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_27),
.B(n_266),
.Y(n_265)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_30),
.A2(n_32),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_30),
.A2(n_161),
.B1(n_163),
.B2(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_30),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_30),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_38),
.A2(n_47),
.B1(n_90),
.B2(n_124),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_40),
.B(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_43),
.A2(n_48),
.B1(n_50),
.B2(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_43),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_43),
.A2(n_50),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_47),
.A2(n_124),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_47),
.A2(n_177),
.B(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_47),
.B(n_156),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_50),
.B(n_178),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_51),
.B(n_64),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_61),
.B2(n_63),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_53),
.B1(n_63),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_52),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_52),
.A2(n_150),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_53),
.A2(n_61),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_53),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_53),
.A2(n_127),
.B(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_SL g157 ( 
.A(n_57),
.B(n_68),
.C(n_74),
.Y(n_157)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_58),
.A2(n_73),
.B(n_155),
.C(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_58),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B(n_77),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_131),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_71),
.A2(n_78),
.B(n_155),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_107),
.B(n_110),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_75),
.A2(n_110),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_83),
.B(n_156),
.CON(n_155),
.SN(n_155)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_96),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B(n_94),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_90),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_90),
.A2(n_227),
.B(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_117)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_130),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_123),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_149),
.B1(n_151),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_166),
.B(n_293),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_164),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_137),
.B(n_164),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_142),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_144),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_152),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_147),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_154),
.B1(n_158),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_156),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_159),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_196),
.B(n_287),
.C(n_292),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_190),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_190),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_180),
.C(n_183),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_169),
.A2(n_170),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_280),
.B(n_286),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_228),
.B(n_279),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_217),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_217),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_210),
.C(n_214),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_202),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_210),
.A2(n_214),
.B1(n_215),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_273),
.B(n_278),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_249),
.B(n_272),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_243),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_277)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_258),
.B(n_271),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_256),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_264),
.B(n_270),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule