module fake_jpeg_14087_n_149 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_30),
.Y(n_32)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_49),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_10),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_27),
.B1(n_12),
.B2(n_29),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_65),
.B1(n_76),
.B2(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_12),
.C(n_29),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_32),
.C(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_62),
.Y(n_95)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_26),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_81),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_30),
.B1(n_16),
.B2(n_3),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.C(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_16),
.B1(n_1),
.B2(n_4),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_84),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_4),
.B1(n_16),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_55),
.B1(n_63),
.B2(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_54),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_88),
.C(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_68),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_56),
.B(n_62),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_106),
.B(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_58),
.C(n_74),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_88),
.C(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_57),
.B1(n_58),
.B2(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_79),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_88),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_97),
.B1(n_110),
.B2(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_109),
.B1(n_107),
.B2(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_117),
.B1(n_120),
.B2(n_115),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_113),
.C(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_98),
.Y(n_134)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_106),
.B1(n_115),
.B2(n_123),
.C(n_127),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_130),
.CI(n_129),
.CON(n_137),
.SN(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_132),
.C(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_141),
.B(n_142),
.Y(n_144)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_140),
.C(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_144),
.C(n_130),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_138),
.B(n_142),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_136),
.Y(n_149)
);


endmodule