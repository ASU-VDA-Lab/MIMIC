module fake_jpeg_28050_n_55 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_SL g22 ( 
.A(n_20),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_22),
.B(n_4),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_22),
.B(n_3),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_2),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_35),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_10),
.B1(n_18),
.B2(n_5),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_8),
.B1(n_16),
.B2(n_6),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_2),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_39),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_7),
.B1(n_11),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_19),
.B1(n_14),
.B2(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_47),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

AO21x1_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_50),
.B(n_49),
.Y(n_55)
);


endmodule