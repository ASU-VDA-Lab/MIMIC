module fake_jpeg_22565_n_26 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_26);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_26;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_17;
wire n_25;
wire n_15;

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

HAxp5_ASAP7_75t_SL g14 ( 
.A(n_0),
.B(n_2),
.CON(n_14),
.SN(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_19),
.C(n_20),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_3),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_22),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_25),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_26)
);


endmodule