module real_jpeg_33335_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_0),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_536),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_1),
.B(n_537),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_4),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_5),
.Y(n_270)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_5),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_251),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_8),
.A2(n_254),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_8),
.A2(n_95),
.B1(n_254),
.B2(n_326),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_8),
.A2(n_254),
.B1(n_436),
.B2(n_438),
.Y(n_435)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

OAI22x1_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_10),
.Y(n_64)
);

AO22x2_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_64),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g231 ( 
.A1(n_10),
.A2(n_64),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_10),
.A2(n_64),
.B1(n_267),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_11),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_12),
.A2(n_29),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_29),
.B1(n_221),
.B2(n_227),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_12),
.A2(n_29),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_13),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_13),
.Y(n_94)
);

AOI22x1_ASAP7_75t_SL g142 ( 
.A1(n_13),
.A2(n_94),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g208 ( 
.A1(n_13),
.A2(n_94),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_13),
.B(n_341),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g400 ( 
.A1(n_13),
.A2(n_401),
.A3(n_407),
.B1(n_409),
.B2(n_413),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_13),
.B(n_140),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_189),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_187),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_175),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_18),
.B(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_149),
.C(n_159),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_20),
.A2(n_149),
.B1(n_174),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_20),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_68),
.Y(n_20)
);

OA21x2_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_35),
.B(n_48),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_22),
.A2(n_150),
.B(n_178),
.Y(n_177)
);

OA21x2_ASAP7_75t_SL g185 ( 
.A1(n_22),
.A2(n_35),
.B(n_48),
.Y(n_185)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_33),
.Y(n_156)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_34),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_34),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_36),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_36),
.B(n_94),
.Y(n_314)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2x1p5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_37),
.B(n_250),
.Y(n_379)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_40),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_42),
.Y(n_355)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_42),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_44),
.Y(n_170)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_49),
.B(n_379),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_50),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_50),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_50),
.A2(n_153),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_50),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_99),
.B(n_148),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_101),
.C(n_138),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_185),
.C(n_186),
.Y(n_184)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_69),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_69),
.B(n_376),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_69),
.B(n_376),
.C(n_378),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_81),
.B(n_91),
.Y(n_69)
);

AO22x2_ASAP7_75t_L g219 ( 
.A1(n_70),
.A2(n_81),
.B1(n_220),
.B2(n_231),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_70),
.B(n_91),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_70),
.B(n_220),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_70),
.B(n_325),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_70),
.B(n_231),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_70),
.Y(n_451)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_82),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_74),
.Y(n_421)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_76),
.Y(n_272)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_76),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_76),
.Y(n_412)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_81),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_81),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_81),
.B(n_91),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_85),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_85),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_90),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_93),
.Y(n_233)
);

OAI21x1_ASAP7_75t_SL g153 ( 
.A1(n_94),
.A2(n_154),
.B(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_158),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g330 ( 
.A1(n_94),
.A2(n_331),
.A3(n_334),
.B1(n_339),
.B2(n_340),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_94),
.B(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_94),
.B(n_451),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_94),
.B(n_199),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_97),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_98),
.Y(n_328)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_137),
.Y(n_99)
);

NAND2x1_ASAP7_75t_L g239 ( 
.A(n_100),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_102),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_140),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_103),
.B(n_140),
.Y(n_276)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_106),
.Y(n_307)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_106),
.Y(n_351)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_111),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_112),
.B(n_142),
.Y(n_275)
);

AO21x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_121),
.B(n_129),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_113),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_116),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_130),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_139),
.B(n_304),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_140),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_140),
.B(n_305),
.Y(n_377)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_171),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_149),
.A2(n_174),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_150),
.B(n_249),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_151),
.B(n_153),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_152),
.B(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_157),
.Y(n_365)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_160),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_173),
.C(n_174),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_162),
.B(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_171),
.B(n_172),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_169),
.A2(n_361),
.B(n_365),
.Y(n_360)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_179),
.B(n_497),
.C(n_498),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_180),
.B(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_296),
.B(n_533),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_290),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_277),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_192),
.B(n_277),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_237),
.C(n_245),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_194),
.B(n_238),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_218),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_195)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g329 ( 
.A(n_196),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_196),
.A2(n_216),
.B1(n_330),
.B2(n_388),
.Y(n_387)
);

AO21x2_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B(n_207),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g485 ( 
.A1(n_197),
.A2(n_318),
.B(n_368),
.Y(n_485)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_198),
.B(n_208),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_198),
.B(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_214),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_216),
.A2(n_219),
.B1(n_279),
.B2(n_510),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_218),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_219),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_242),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_243),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_243),
.B(n_261),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_244),
.B(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_246),
.B(n_514),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_259),
.C(n_273),
.Y(n_246)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_248),
.B(n_274),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_260),
.B(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_262),
.B(n_493),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_263),
.B(n_434),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_265),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_265),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_270),
.Y(n_370)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2x1p5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_275),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_276),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_288),
.C(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_290),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

NOR2x1_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_291),
.B(n_293),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_523),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_471),
.B(n_522),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_380),
.B(n_470),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_343),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_300),
.B(n_343),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_323),
.C(n_329),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_301),
.A2(n_302),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_313),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_322),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_312),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B(n_322),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_315),
.Y(n_346)
);

NOR2x1p5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_316),
.Y(n_455)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_318),
.B(n_434),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_319),
.Y(n_367)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_329),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_324),
.B(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_374),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_345),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_347),
.B(n_374),
.C(n_501),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_366),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_348),
.B(n_366),
.Y(n_477)
);

OAI31xp33_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_352),
.A3(n_356),
.B(n_360),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_391),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_395),
.B(n_469),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_382),
.B(n_385),
.Y(n_469)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.C(n_392),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_387),
.B(n_465),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_389),
.A2(n_390),
.B1(n_392),
.B2(n_393),
.Y(n_465)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_424),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_463),
.B(n_468),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_441),
.B(n_462),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_425),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_425),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_422),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_400),
.B1(n_422),
.B2(n_423),
.Y(n_447)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_424),
.B(n_431),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_432),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_433),
.C(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_448),
.B(n_461),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_447),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_447),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_455),
.Y(n_454)
);

BUFx4f_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_453),
.B(n_460),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_452),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_466),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_504),
.C(n_515),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_499),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_487),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_474),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_483),
.C(n_484),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_482),
.C(n_491),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

XOR2x1_ASAP7_75t_SL g503 ( 
.A(n_483),
.B(n_484),
.Y(n_503)
);

XOR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_486),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_494),
.B2(n_495),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_490),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_517),
.C(n_519),
.Y(n_516)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_502),
.Y(n_526)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_513),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_505),
.B(n_513),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_509),
.C(n_511),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_509),
.Y(n_521)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_521),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_515),
.A2(n_525),
.B(n_527),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_520),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_520),
.Y(n_531)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_530),
.B(n_532),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);


endmodule