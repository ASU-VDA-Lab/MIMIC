module fake_jpeg_8880_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_13),
.B1(n_9),
.B2(n_16),
.Y(n_31)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_12),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_12),
.C(n_9),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_31),
.B(n_22),
.C(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_48),
.B1(n_32),
.B2(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

XOR2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_53),
.B(n_58),
.Y(n_69)
);

XOR2x1_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_60),
.B1(n_27),
.B2(n_28),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_50),
.C(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_47),
.B(n_42),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_65),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_57),
.A3(n_61),
.B1(n_55),
.B2(n_41),
.C(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_15),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_27),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_28),
.C(n_17),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_10),
.C(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_76),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_62),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_80),
.C(n_0),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_63),
.B1(n_68),
.B2(n_15),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_10),
.B(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_83),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_75),
.B(n_70),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_75),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_39),
.C1(n_76),
.C2(n_79),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_90),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_89),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_7),
.Y(n_93)
);


endmodule