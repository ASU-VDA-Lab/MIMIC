module fake_jpeg_13019_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AND2x6_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_40),
.B(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_37),
.Y(n_92)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_1),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_32),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_21),
.B1(n_32),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_75),
.B1(n_52),
.B2(n_3),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_61),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_30),
.B1(n_38),
.B2(n_34),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_80),
.B1(n_64),
.B2(n_19),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_39),
.B1(n_38),
.B2(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_39),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_34),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_37),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_61),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_53),
.B1(n_50),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_68),
.B1(n_86),
.B2(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_21),
.B1(n_22),
.B2(n_56),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_129),
.B1(n_106),
.B2(n_101),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_119),
.Y(n_148)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_121),
.Y(n_156)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_125),
.Y(n_143)
);

BUFx2_ASAP7_75t_SL g125 ( 
.A(n_69),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_52),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_1),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_5),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_100),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_2),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_75),
.B1(n_96),
.B2(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_118),
.B1(n_110),
.B2(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_103),
.A2(n_89),
.B1(n_82),
.B2(n_70),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_142),
.B1(n_149),
.B2(n_9),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_82),
.B1(n_70),
.B2(n_95),
.Y(n_142)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_67),
.A3(n_86),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_7),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_150),
.B(n_151),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_2),
.C(n_3),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_95),
.C(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_5),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_8),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_161),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_141),
.B1(n_140),
.B2(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_117),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_123),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_167),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_111),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_114),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_136),
.B1(n_153),
.B2(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_137),
.B(n_139),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_146),
.C(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_181),
.C(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_169),
.B(n_157),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_135),
.C(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NOR2x1_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_168),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_151),
.C(n_152),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_198),
.B1(n_182),
.B2(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_167),
.C(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_206),
.C(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

OA21x2_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_207),
.B(n_147),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_172),
.C(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_180),
.A3(n_188),
.B1(n_185),
.B2(n_193),
.C1(n_182),
.C2(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

AOI321xp33_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_190),
.A3(n_179),
.B1(n_175),
.B2(n_194),
.C(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_199),
.B1(n_191),
.B2(n_203),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_175),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_225),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_216),
.C(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_195),
.C(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_174),
.B1(n_160),
.B2(n_187),
.Y(n_225)
);

AOI31xp67_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_212),
.A3(n_214),
.B(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_227),
.B1(n_162),
.B2(n_166),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_230),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_209),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_165),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_215),
.B(n_219),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_235),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_233),
.A2(n_230),
.B(n_166),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_9),
.B(n_155),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.C(n_236),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_155),
.Y(n_242)
);


endmodule