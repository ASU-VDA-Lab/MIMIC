module fake_jpeg_26030_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_31),
.Y(n_59)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_36),
.B1(n_41),
.B2(n_37),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_69),
.B1(n_28),
.B2(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_59),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_28),
.B(n_5),
.Y(n_100)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_32),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_28),
.B(n_16),
.C(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_65),
.B1(n_28),
.B2(n_16),
.Y(n_86)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_34),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_24),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_48),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_43),
.Y(n_77)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_79),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_81),
.B(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_93),
.B1(n_71),
.B2(n_66),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_14),
.C(n_13),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_27),
.B1(n_28),
.B2(n_16),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_64),
.B1(n_72),
.B2(n_61),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_43),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_71),
.C(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_95),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_2),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_102),
.B(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_3),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_3),
.B(n_6),
.C(n_7),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_120),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_117),
.B1(n_125),
.B2(n_127),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_85),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_61),
.B1(n_60),
.B2(n_64),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_124),
.C(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_71),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_102),
.B(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_54),
.C(n_51),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_54),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_75),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_54),
.B1(n_66),
.B2(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_76),
.A2(n_66),
.B1(n_8),
.B2(n_11),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_103),
.B1(n_83),
.B2(n_11),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_82),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_75),
.B1(n_84),
.B2(n_80),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_107),
.B1(n_128),
.B2(n_122),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_146),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_93),
.Y(n_142)
);

XOR2x1_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_91),
.C(n_73),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_150),
.C(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_97),
.C(n_73),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_112),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_83),
.B1(n_111),
.B2(n_130),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_161),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_152),
.B(n_148),
.C(n_150),
.D(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_173),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_142),
.B(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_110),
.B1(n_107),
.B2(n_104),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_110),
.B1(n_107),
.B2(n_104),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_159),
.A3(n_171),
.B1(n_164),
.B2(n_158),
.C1(n_134),
.C2(n_166),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_127),
.B1(n_113),
.B2(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_144),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_143),
.B(n_155),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_170),
.CI(n_163),
.CON(n_189),
.SN(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_181),
.C(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.C(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_167),
.C(n_149),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_161),
.B1(n_160),
.B2(n_147),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_200),
.B1(n_191),
.B2(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_205),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_177),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_180),
.A3(n_182),
.B1(n_188),
.B2(n_94),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_208),
.B1(n_197),
.B2(n_189),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_7),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_198),
.C(n_199),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_7),
.B(n_8),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_11),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_194),
.C(n_190),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_193),
.C(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_213),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_203),
.B1(n_208),
.B2(n_209),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_196),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_212),
.Y(n_222)
);

OAI221xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_197),
.B1(n_207),
.B2(n_196),
.C(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_218),
.B(n_210),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_213),
.B(n_216),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_12),
.Y(n_227)
);


endmodule