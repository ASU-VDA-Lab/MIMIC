module fake_jpeg_4820_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_28),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_62),
.B1(n_29),
.B2(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_41),
.B1(n_17),
.B2(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_94),
.B1(n_35),
.B2(n_23),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_36),
.B(n_44),
.C(n_16),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_43),
.B1(n_36),
.B2(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_84),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_36),
.B1(n_44),
.B2(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_90),
.B1(n_24),
.B2(n_21),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_50),
.Y(n_108)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_91),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_16),
.B1(n_45),
.B2(n_18),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_92),
.B1(n_22),
.B2(n_21),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_21),
.B1(n_22),
.B2(n_34),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_19),
.B1(n_23),
.B2(n_35),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_24),
.B1(n_31),
.B2(n_34),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_18),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_104),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_130),
.B1(n_72),
.B2(n_70),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_37),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_51),
.B1(n_19),
.B2(n_27),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_94),
.B1(n_79),
.B2(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_45),
.B1(n_46),
.B2(n_39),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_71),
.B1(n_18),
.B2(n_39),
.Y(n_131)
);

AO21x2_ASAP7_75t_SL g192 ( 
.A1(n_131),
.A2(n_39),
.B(n_46),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_42),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_143),
.C(n_108),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_37),
.C(n_38),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_151),
.B1(n_104),
.B2(n_121),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_26),
.B(n_102),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_81),
.B1(n_98),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_159),
.B1(n_112),
.B2(n_121),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_37),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_107),
.B1(n_104),
.B2(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_174),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_146),
.A3(n_137),
.B1(n_134),
.B2(n_149),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_187),
.C(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_112),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_102),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_37),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_182),
.B2(n_194),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_177),
.A2(n_25),
.B1(n_33),
.B2(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_186),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_115),
.B(n_101),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_193),
.B1(n_158),
.B2(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_130),
.B1(n_127),
.B2(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2x1p5_ASAP7_75t_SL g185 ( 
.A(n_131),
.B(n_33),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_192),
.B(n_82),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_137),
.A2(n_134),
.B(n_154),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_114),
.C(n_113),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_135),
.A2(n_86),
.B(n_116),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_159),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_114),
.C(n_116),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_140),
.A2(n_123),
.B1(n_105),
.B2(n_46),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_123),
.B1(n_105),
.B2(n_67),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_204),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_201),
.B(n_210),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_192),
.B1(n_181),
.B2(n_162),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_203),
.A2(n_222),
.B1(n_165),
.B2(n_174),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_217),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_145),
.B1(n_93),
.B2(n_160),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_224),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_38),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_142),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_218),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_161),
.B(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_187),
.C(n_191),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_75),
.B(n_38),
.C(n_37),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_189),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_87),
.A3(n_33),
.B1(n_25),
.B2(n_10),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_176),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_33),
.B1(n_87),
.B2(n_2),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_186),
.B(n_190),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_234),
.B1(n_196),
.B2(n_207),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_235),
.B1(n_237),
.B2(n_206),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_218),
.B(n_202),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_180),
.B1(n_188),
.B2(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_203),
.B1(n_222),
.B2(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_170),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_246),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_244),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_173),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_252),
.A2(n_256),
.B(n_5),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_241),
.B(n_251),
.Y(n_283)
);

AOI21x1_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_215),
.B(n_209),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_217),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_258),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_216),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_197),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_239),
.CI(n_227),
.CON(n_275),
.SN(n_275)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_216),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_263),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_237),
.B(n_215),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_195),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_15),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_1),
.C(n_3),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_3),
.C(n_5),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_244),
.B1(n_12),
.B2(n_10),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_15),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_5),
.C(n_6),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_233),
.C(n_6),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_234),
.B(n_248),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_227),
.B(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_250),
.B1(n_241),
.B2(n_238),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_289),
.B1(n_269),
.B2(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_290),
.C(n_268),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_228),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_228),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_13),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_7),
.C(n_8),
.Y(n_290)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_293),
.B(n_277),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_255),
.B1(n_258),
.B2(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_275),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_255),
.C(n_266),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_299),
.C(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_254),
.C(n_8),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_8),
.C(n_12),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_8),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_304),
.CI(n_287),
.CON(n_310),
.SN(n_310)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_13),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_273),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_308),
.C(n_311),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_288),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B(n_316),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_290),
.C(n_277),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_315),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_273),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_274),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_281),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_295),
.B(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_302),
.B1(n_292),
.B2(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_322),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_293),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_308),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_291),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_325),
.B(n_283),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_306),
.A2(n_289),
.B(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_318),
.B(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_330),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_332),
.B1(n_326),
.B2(n_323),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_313),
.B(n_329),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_334),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_333),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_284),
.B(n_13),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_14),
.B1(n_204),
.B2(n_302),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_340),
.Y(n_341)
);


endmodule