module real_jpeg_30167_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_285, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_285;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_283;
wire n_85;
wire n_81;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_273;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_0),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_4),
.B1(n_18),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_22),
.B1(n_25),
.B2(n_43),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_22),
.B(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_43),
.B1(n_69),
.B2(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_21),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_5),
.B(n_49),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_66),
.B(n_70),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_48),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_4),
.A2(n_10),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_4),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_9),
.B1(n_18),
.B2(n_32),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_8),
.B1(n_18),
.B2(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_23),
.B(n_43),
.C(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_22),
.B1(n_25),
.B2(n_50),
.Y(n_53)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_58),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_9),
.A2(n_32),
.B1(n_49),
.B2(n_51),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_17),
.B1(n_49),
.B2(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_10),
.A2(n_17),
.B1(n_69),
.B2(n_70),
.Y(n_208)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_11),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_35),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_33),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_28),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_21),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_20),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_21),
.A2(n_26),
.B1(n_42),
.B2(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_22),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_22),
.A2(n_43),
.B(n_146),
.C(n_147),
.Y(n_145)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_29),
.B(n_37),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_40),
.B(n_41),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_73),
.B(n_283),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_38),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_38),
.B(n_281),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_44),
.CI(n_54),
.CON(n_38),
.SN(n_38)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_41),
.B(n_57),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_42),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_43),
.A2(n_49),
.B(n_67),
.C(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_43),
.B(n_100),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_43),
.B(n_68),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_47),
.B(n_85),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_48),
.A2(n_60),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_51),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_86),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_61),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_55),
.B(n_89),
.C(n_90),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_55),
.A2(n_88),
.B1(n_104),
.B2(n_129),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_55),
.B(n_129),
.C(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_55),
.A2(n_88),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_59),
.A2(n_61),
.B1(n_262),
.B2(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_59),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_61),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_61),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_64),
.A2(n_68),
.B1(n_109),
.B2(n_116),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_64),
.A2(n_68),
.B1(n_72),
.B2(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_68),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_69),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_97),
.Y(n_96)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_280),
.B(n_282),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_254),
.A3(n_273),
.B1(n_278),
.B2(n_279),
.C(n_285),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_237),
.B(n_253),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_218),
.B(n_236),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_139),
.B(n_201),
.C(n_217),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_126),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_79),
.B(n_126),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_101),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_80),
.B(n_102),
.C(n_112),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_136),
.C(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_89),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_82),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_82),
.B(n_243),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_87),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_94),
.A2(n_134),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_94),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_94),
.B(n_184),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_94),
.B(n_161),
.C(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_97),
.B(n_123),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_97),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_96),
.A2(n_100),
.B1(n_121),
.B2(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_111),
.B2(n_112),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_129),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_105),
.Y(n_261)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_110),
.A2(n_130),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_110),
.A2(n_130),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_110),
.A2(n_130),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_110),
.B(n_260),
.C(n_262),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_110),
.B(n_267),
.C(n_272),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_113),
.A2(n_114),
.B1(n_168),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_113),
.B(n_120),
.Y(n_211)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_129),
.C(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_114),
.B(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B(n_118),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_118),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_135),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_211),
.C(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_135),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_136),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_200),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_194),
.B(n_199),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_164),
.B(n_193),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_152),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_151),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_158),
.B2(n_159),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_161),
.C(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_155),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_156),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_163),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_163),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_207),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_188),
.B(n_192),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_175),
.B(n_187),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_170),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B(n_186),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_185),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_216),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_210),
.C(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_220),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_227),
.C(n_235),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_232),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_246),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_239),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_251),
.B2(n_252),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_245),
.C(n_252),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_256),
.C(n_263),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_256),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_265),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_264),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);


endmodule