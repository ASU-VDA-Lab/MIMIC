module fake_jpeg_16199_n_351 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_76),
.B1(n_29),
.B2(n_28),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_21),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_70),
.B(n_29),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_74),
.B1(n_29),
.B2(n_28),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_32),
.B1(n_24),
.B2(n_31),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_98),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_106),
.B1(n_73),
.B2(n_62),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_63),
.B(n_25),
.Y(n_134)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_79),
.B1(n_80),
.B2(n_54),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_108),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_33),
.B1(n_53),
.B2(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_26),
.C(n_14),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_53),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_24),
.B(n_31),
.C(n_30),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_111),
.Y(n_142)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_42),
.B1(n_24),
.B2(n_30),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_33),
.B1(n_74),
.B2(n_27),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_70),
.C(n_51),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_138),
.C(n_20),
.Y(n_154)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_128),
.B1(n_136),
.B2(n_100),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_73),
.B1(n_66),
.B2(n_59),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_132),
.B1(n_137),
.B2(n_104),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_25),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_133),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_54),
.B1(n_80),
.B2(n_59),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_56),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_141),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_65),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_82),
.B1(n_90),
.B2(n_93),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_37),
.A3(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_33),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_91),
.B1(n_109),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_155),
.B1(n_167),
.B2(n_113),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_156),
.B1(n_168),
.B2(n_165),
.Y(n_171)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_161),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_116),
.Y(n_192)
);

XNOR2x2_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_84),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_132),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_165),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_168),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_93),
.C(n_19),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_113),
.B1(n_117),
.B2(n_128),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_35),
.C(n_22),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_35),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_35),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_110),
.B1(n_103),
.B2(n_95),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_157),
.B(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_95),
.B1(n_11),
.B2(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_35),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_134),
.B1(n_140),
.B2(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_173),
.B(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_179),
.B1(n_184),
.B2(n_37),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_125),
.B1(n_123),
.B2(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_129),
.B1(n_135),
.B2(n_130),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_191),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_147),
.B1(n_167),
.B2(n_160),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_113),
.B1(n_124),
.B2(n_117),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_19),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.C(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_158),
.B(n_149),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_127),
.B(n_1),
.Y(n_193)
);

AND2x4_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_116),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_145),
.B1(n_144),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_145),
.B1(n_127),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_203),
.B1(n_206),
.B2(n_213),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_212),
.C(n_220),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_153),
.B1(n_124),
.B2(n_151),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_169),
.B1(n_83),
.B2(n_120),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_209),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_126),
.B1(n_122),
.B2(n_37),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_126),
.C(n_122),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_35),
.B1(n_22),
.B2(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_35),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_175),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_35),
.B1(n_23),
.B2(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_23),
.C(n_9),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_227),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_172),
.C(n_188),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_238),
.C(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_190),
.C(n_179),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_180),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_219),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_187),
.B(n_193),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_216),
.B(n_214),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_211),
.B1(n_197),
.B2(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_247),
.C(n_230),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_196),
.C(n_218),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_264),
.C(n_231),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_211),
.B1(n_203),
.B2(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_206),
.B1(n_217),
.B2(n_198),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_213),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_220),
.B1(n_175),
.B2(n_185),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_230),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_23),
.C(n_3),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_224),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_274),
.C(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_225),
.C(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_262),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_233),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_225),
.C(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_286),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_232),
.C(n_228),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_284),
.C(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_228),
.C(n_226),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_245),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_226),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_266),
.B1(n_260),
.B2(n_245),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_266),
.B1(n_251),
.B2(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_291),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_297),
.C(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_253),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_249),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_263),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_269),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_23),
.C(n_6),
.Y(n_314)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_307),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_271),
.B1(n_280),
.B2(n_268),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_309),
.B1(n_293),
.B2(n_13),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_251),
.B1(n_260),
.B2(n_282),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_282),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_5),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_23),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_297),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_294),
.B1(n_290),
.B2(n_302),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_326),
.B1(n_315),
.B2(n_303),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_327),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_293),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_323),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_6),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_316),
.C(n_307),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_306),
.A2(n_9),
.B(n_10),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_335),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_334),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_308),
.C(n_16),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_6),
.C(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_329),
.B(n_336),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_338),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_332),
.A2(n_320),
.B(n_325),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_340),
.A2(n_7),
.B(n_8),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_323),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_345),
.B(n_346),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_341),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_342),
.C(n_339),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_7),
.B(n_8),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_8),
.Y(n_351)
);


endmodule