module fake_jpeg_10760_n_433 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_433);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_20),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_63),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g128 ( 
.A(n_67),
.Y(n_128)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_31),
.B1(n_23),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_86),
.A2(n_139),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_42),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_103),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_28),
.B1(n_27),
.B2(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_90),
.A2(n_100),
.B1(n_125),
.B2(n_86),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_30),
.B1(n_25),
.B2(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_42),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_39),
.B(n_19),
.C(n_32),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_16),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_21),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_53),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_45),
.B(n_34),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_58),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_39),
.B(n_32),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_21),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_37),
.C(n_19),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_29),
.Y(n_123)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_28),
.B1(n_25),
.B2(n_30),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_38),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_36),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_80),
.B(n_28),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_12),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_47),
.A2(n_37),
.B1(n_35),
.B2(n_25),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_45),
.Y(n_140)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_94),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_R g237 ( 
.A(n_147),
.B(n_195),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_153),
.B1(n_154),
.B2(n_162),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_151),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_35),
.B1(n_18),
.B2(n_24),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_35),
.B1(n_18),
.B2(n_24),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_174),
.Y(n_230)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_40),
.B1(n_24),
.B2(n_22),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_118),
.B1(n_122),
.B2(n_90),
.Y(n_162)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_120),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_40),
.B1(n_22),
.B2(n_35),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_132),
.B1(n_115),
.B2(n_104),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_40),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_182),
.C(n_107),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_172),
.B(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_0),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_0),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_115),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_180),
.B1(n_198),
.B2(n_102),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_1),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_185),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_187),
.B(n_191),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_83),
.Y(n_199)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_12),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_98),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_107),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_87),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_199),
.B(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_218),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_128),
.CI(n_127),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_203),
.B(n_232),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_102),
.B1(n_108),
.B2(n_112),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_205),
.A2(n_227),
.B1(n_228),
.B2(n_246),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_142),
.B(n_93),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_114),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_93),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_211),
.B(n_245),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_225),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_112),
.B1(n_124),
.B2(n_95),
.Y(n_213)
);

OR2x6_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_124),
.Y(n_216)
);

NAND2x1p5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_182),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_150),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_149),
.A2(n_91),
.B1(n_134),
.B2(n_11),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_171),
.A2(n_172),
.B1(n_195),
.B2(n_163),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_161),
.A2(n_91),
.B1(n_134),
.B2(n_127),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_163),
.B(n_134),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_142),
.B(n_127),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_235),
.A2(n_212),
.B1(n_216),
.B2(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_161),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_163),
.B1(n_143),
.B2(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_181),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_159),
.B(n_173),
.C(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_181),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_247),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_145),
.B(n_157),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_168),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_165),
.B(n_184),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_182),
.B(n_178),
.C(n_187),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_211),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_252),
.B(n_255),
.Y(n_300)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_258),
.B(n_216),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_210),
.A2(n_144),
.B(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_169),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_263),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_201),
.A2(n_189),
.B1(n_177),
.B2(n_191),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_266),
.A2(n_268),
.B1(n_282),
.B2(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_201),
.A2(n_192),
.B1(n_146),
.B2(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_241),
.B(n_146),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_275),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_167),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_221),
.A2(n_185),
.B1(n_156),
.B2(n_158),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_227),
.B1(n_223),
.B2(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_285),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_209),
.A2(n_216),
.B1(n_221),
.B2(n_239),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_222),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_206),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_204),
.B(n_236),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_240),
.B(n_238),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_290),
.B(n_274),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_204),
.B(n_215),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_203),
.B(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_219),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_229),
.C(n_240),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_324),
.C(n_327),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_216),
.B1(n_228),
.B2(n_203),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_310),
.B1(n_311),
.B2(n_287),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_309),
.B1(n_314),
.B2(n_285),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_256),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_305),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_276),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g351 ( 
.A1(n_303),
.A2(n_312),
.B(n_307),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_261),
.A2(n_237),
.B(n_205),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_283),
.B1(n_266),
.B2(n_268),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_279),
.A2(n_237),
.B1(n_235),
.B2(n_214),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_281),
.A2(n_223),
.B1(n_217),
.B2(n_206),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_223),
.B(n_217),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_313),
.B(n_303),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_261),
.A2(n_284),
.B1(n_264),
.B2(n_280),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_250),
.A2(n_276),
.B1(n_290),
.B2(n_292),
.Y(n_314)
);

A2O1A1O1Ixp25_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_291),
.B(n_267),
.C(n_288),
.D(n_257),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_276),
.C(n_273),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_267),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_334),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_306),
.B(n_251),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_332),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_333),
.B1(n_354),
.B2(n_348),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_296),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_308),
.A2(n_257),
.B1(n_272),
.B2(n_255),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_334),
.B(n_315),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_335),
.A2(n_341),
.B1(n_343),
.B2(n_353),
.Y(n_365)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_262),
.B1(n_265),
.B2(n_269),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_319),
.B1(n_315),
.B2(n_322),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_253),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_346),
.C(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_321),
.A2(n_310),
.B1(n_294),
.B2(n_305),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_259),
.B1(n_277),
.B2(n_254),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_286),
.C(n_270),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_293),
.C(n_299),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_321),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_349),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_301),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_300),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_304),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_351),
.A2(n_352),
.B(n_355),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_308),
.B1(n_309),
.B2(n_325),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_320),
.A2(n_301),
.B1(n_298),
.B2(n_326),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_296),
.A2(n_319),
.B(n_317),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g356 ( 
.A1(n_330),
.A2(n_304),
.B1(n_317),
.B2(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_364),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_362),
.A2(n_367),
.B1(n_360),
.B2(n_359),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_352),
.A2(n_322),
.B(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_353),
.A2(n_341),
.B1(n_335),
.B2(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_371),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_328),
.A2(n_349),
.B(n_342),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_372),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_350),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_373),
.B(n_375),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_374),
.C(n_361),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_358),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_380),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_375),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_347),
.B1(n_338),
.B2(n_339),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_391),
.B1(n_395),
.B2(n_376),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_368),
.B(n_338),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_372),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_356),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_377),
.C(n_364),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_365),
.C(n_366),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_371),
.A2(n_363),
.B1(n_370),
.B2(n_365),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_356),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_387),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_379),
.B(n_381),
.Y(n_397)
);

AOI21x1_ASAP7_75t_SL g415 ( 
.A1(n_397),
.A2(n_407),
.B(n_382),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_369),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_402),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_399),
.B(n_400),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_357),
.C(n_359),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_383),
.C(n_390),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_357),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_380),
.A2(n_360),
.B1(n_376),
.B2(n_379),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_409),
.B1(n_389),
.B2(n_398),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_406),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_381),
.B1(n_393),
.B2(n_386),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_391),
.A2(n_395),
.B1(n_393),
.B2(n_387),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_396),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_403),
.B1(n_400),
.B2(n_397),
.Y(n_419)
);

AOI21xp33_ASAP7_75t_L g413 ( 
.A1(n_404),
.A2(n_385),
.B(n_382),
.Y(n_413)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_413),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_420),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_399),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_401),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_423),
.B(n_411),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_425),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_408),
.C(n_405),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_426),
.A2(n_421),
.B(n_422),
.Y(n_428)
);

NAND4xp25_ASAP7_75t_SL g429 ( 
.A(n_428),
.B(n_410),
.C(n_415),
.D(n_412),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_408),
.B(n_410),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_SL g431 ( 
.A1(n_430),
.A2(n_422),
.B(n_420),
.C(n_427),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_416),
.B(n_409),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_417),
.Y(n_433)
);


endmodule