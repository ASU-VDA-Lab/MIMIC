module fake_jpeg_7744_n_299 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_41),
.B1(n_31),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_62),
.B1(n_53),
.B2(n_47),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_31),
.B1(n_33),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_58),
.B1(n_65),
.B2(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_61),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_64),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_59),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_33),
.C(n_21),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_32),
.C(n_22),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_31),
.B1(n_20),
.B2(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_24),
.B1(n_16),
.B2(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_34),
.B(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_27),
.B(n_29),
.C(n_22),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_77),
.B1(n_46),
.B2(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_9),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_54),
.B(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_82),
.B1(n_91),
.B2(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_52),
.B1(n_46),
.B2(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_44),
.B1(n_19),
.B2(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_54),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_78),
.CI(n_75),
.CON(n_102),
.SN(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_109),
.B(n_19),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_11),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_76),
.B(n_88),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_63),
.B1(n_44),
.B2(n_17),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_68),
.B1(n_79),
.B2(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_55),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_30),
.B(n_28),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_121),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_85),
.B(n_91),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_127),
.B(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_123),
.B1(n_141),
.B2(n_142),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_135),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_71),
.B(n_30),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_107),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_13),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_105),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_30),
.B1(n_50),
.B2(n_26),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_25),
.Y(n_167)
);

CKINVDCx12_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_102),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.C(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_101),
.C(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_108),
.B1(n_102),
.B2(n_98),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_154),
.B1(n_159),
.B2(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_106),
.B1(n_111),
.B2(n_94),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_124),
.B1(n_120),
.B2(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_106),
.B1(n_94),
.B2(n_90),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_128),
.B(n_123),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_30),
.B(n_28),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_165),
.B(n_142),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_28),
.B(n_18),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_28),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_28),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_25),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_141),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_182),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_189),
.Y(n_206)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_179),
.Y(n_210)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_164),
.B(n_160),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_144),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_143),
.C(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_159),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_126),
.CI(n_143),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_184),
.B(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_127),
.B1(n_143),
.B2(n_128),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_192),
.B1(n_196),
.B2(n_165),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_166),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_126),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_125),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_127),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_197),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_125),
.C(n_138),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_200),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_147),
.B1(n_158),
.B2(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_212),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_220),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_153),
.B1(n_158),
.B2(n_155),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_204),
.B1(n_219),
.B2(n_18),
.Y(n_230)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_18),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_171),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_218),
.B1(n_197),
.B2(n_183),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_166),
.B1(n_142),
.B2(n_19),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_142),
.B1(n_1),
.B2(n_0),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_142),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_175),
.C(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_224),
.C(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_175),
.C(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_18),
.C(n_1),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_8),
.B1(n_15),
.B2(n_2),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_239),
.B1(n_201),
.B2(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_18),
.C(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_9),
.C(n_3),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_236),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_0),
.C(n_3),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_208),
.B(n_211),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_250),
.B(n_233),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_237),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_210),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_222),
.C(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_203),
.B1(n_207),
.B2(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_253),
.Y(n_256)
);

OAI22x1_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_205),
.B1(n_200),
.B2(n_220),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_198),
.B1(n_213),
.B2(n_219),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_236),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.C(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_231),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_244),
.B(n_247),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_5),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_7),
.C(n_8),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_274),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_248),
.B1(n_243),
.B2(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_264),
.B(n_10),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_247),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_242),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_260),
.Y(n_282)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_7),
.C(n_10),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_269),
.C(n_11),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_275),
.B1(n_270),
.B2(n_278),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_270),
.B1(n_277),
.B2(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.C(n_292),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_10),
.B(n_11),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_12),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_289),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_295),
.B1(n_290),
.B2(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_279),
.C(n_14),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_279),
.Y(n_299)
);


endmodule