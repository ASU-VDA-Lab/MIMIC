module real_jpeg_12300_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_336, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_336;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_30),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_3),
.B(n_21),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_23),
.B(n_85),
.C(n_229),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_155),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_3),
.B(n_53),
.C(n_66),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_3),
.B(n_86),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_3),
.A2(n_121),
.B(n_254),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_155),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_161),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_161),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_161),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_6),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_78),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_78),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_78),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_9),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_88),
.Y(n_175)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_11),
.B(n_24),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_33),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_13),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_130),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_130),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_14),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_74),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_15),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_120)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_32),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_21),
.A2(n_27),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_21),
.A2(n_27),
.B1(n_36),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_22),
.A2(n_73),
.B(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_22),
.A2(n_28),
.B1(n_73),
.B2(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_22),
.B(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_22),
.A2(n_28),
.B1(n_106),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_22),
.A2(n_75),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_22),
.A2(n_28),
.B1(n_129),
.B2(n_200),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_23),
.A2(n_24),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_23),
.A2(n_26),
.A3(n_31),
.B1(n_157),
.B2(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_27),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_28),
.A2(n_129),
.B(n_131),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_28),
.A2(n_31),
.B(n_155),
.C(n_156),
.Y(n_154)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_34),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_35),
.B(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_329),
.B(n_331),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_317),
.B(n_328),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_146),
.B(n_314),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_133),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_108),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_45),
.B(n_108),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_45),
.Y(n_335)
);

FAx1_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_79),
.CI(n_94),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_46),
.B(n_79),
.C(n_94),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_72),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_47),
.A2(n_48),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_51),
.A2(n_55),
.B1(n_120),
.B2(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_51),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_51),
.A2(n_55),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_53),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_52),
.B(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_55),
.B(n_232),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_69),
.B2(n_71),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_64),
.B1(n_71),
.B2(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_63),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_62),
.B(n_244),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_84),
.B(n_155),
.Y(n_229)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_71),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_64),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_64),
.A2(n_71),
.B1(n_125),
.B2(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_64),
.A2(n_71),
.B1(n_224),
.B2(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_70),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_68),
.A2(n_164),
.B(n_166),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_68),
.A2(n_166),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_68),
.B(n_155),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_71),
.B(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_80),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_81),
.A2(n_89),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_81),
.A2(n_89),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_81),
.A2(n_162),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_81),
.A2(n_198),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_86),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_82),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_82),
.A2(n_86),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_86),
.B(n_181),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_89),
.A2(n_160),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_89),
.A2(n_127),
.B(n_180),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_92),
.A2(n_223),
.B(n_225),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_92),
.A2(n_225),
.B(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_101),
.C(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_101),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_101),
.B(n_138),
.C(n_142),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_105),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_105),
.B(n_137),
.C(n_144),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_115),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_114),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_115),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.C(n_128),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_116),
.A2(n_117),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_122),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_121),
.A2(n_122),
.B1(n_175),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_121),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_122),
.A2(n_185),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_122),
.A2(n_231),
.B(n_259),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_122),
.B(n_155),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_126),
.B(n_128),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_154),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_133),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_145),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_134),
.B(n_145),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_139),
.Y(n_323)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_308),
.B(n_313),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_296),
.B(n_307),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_203),
.A3(n_215),
.B1(n_294),
.B2(n_295),
.C(n_336),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_186),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_150),
.B(n_186),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_169),
.C(n_178),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_151),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_168),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_159),
.C(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_178),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_204),
.B(n_205),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_214),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_207),
.B(n_209),
.C(n_214),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_235),
.B(n_293),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_233),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_217),
.B(n_233),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_218),
.A2(n_219),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_228),
.B(n_230),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_286),
.B(n_292),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_274),
.B(n_285),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_255),
.B(n_273),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_250),
.C(n_252),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_251),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_263),
.B(n_272),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_261),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_267),
.B(n_271),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_281),
.C(n_284),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_306),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_306),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_327),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);


endmodule