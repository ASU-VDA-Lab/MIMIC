module real_aes_10977_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g991 ( .A(n_0), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_0), .A2(n_248), .B1(n_671), .B2(n_1020), .Y(n_1019) );
AO221x1_ASAP7_75t_L g1124 ( .A1(n_1), .A2(n_147), .B1(n_1095), .B2(n_1125), .C(n_1127), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_2), .A2(n_224), .B1(n_327), .B2(n_328), .Y(n_326) );
INVxp33_ASAP7_75t_L g378 ( .A(n_2), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_3), .A2(n_99), .B1(n_603), .B2(n_1403), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_3), .A2(n_99), .B1(n_677), .B2(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g462 ( .A(n_4), .Y(n_462) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_5), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_5), .A2(n_209), .B1(n_671), .B2(n_867), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_6), .A2(n_172), .B1(n_475), .B2(n_573), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_6), .A2(n_126), .B1(n_401), .B2(n_440), .C(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_7), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_7), .B(n_195), .Y(n_283) );
AND2x2_ASAP7_75t_L g387 ( .A(n_7), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g461 ( .A(n_7), .Y(n_461) );
INVx1_ASAP7_75t_L g699 ( .A(n_8), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_8), .A2(n_185), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_9), .A2(n_15), .B1(n_500), .B2(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g538 ( .A(n_9), .Y(n_538) );
OA22x2_ASAP7_75t_L g614 ( .A1(n_10), .A2(n_615), .B1(n_689), .B2(n_690), .Y(n_614) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_10), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_10), .A2(n_105), .B1(n_1095), .B2(n_1099), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_11), .A2(n_47), .B1(n_439), .B2(n_717), .Y(n_721) );
INVx1_ASAP7_75t_L g759 ( .A(n_11), .Y(n_759) );
INVxp67_ASAP7_75t_L g999 ( .A(n_12), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_12), .A2(n_75), .B1(n_652), .B2(n_671), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_13), .A2(n_95), .B1(n_328), .B2(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g598 ( .A(n_13), .Y(n_598) );
OAI332xp33_ASAP7_75t_L g626 ( .A1(n_14), .A2(n_420), .A3(n_457), .B1(n_627), .B2(n_631), .B3(n_636), .C1(n_643), .C2(n_648), .Y(n_626) );
INVx1_ASAP7_75t_L g685 ( .A(n_14), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_15), .A2(n_108), .B1(n_533), .B2(n_535), .C(n_537), .Y(n_532) );
INVxp67_ASAP7_75t_L g888 ( .A(n_16), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g916 ( .A1(n_16), .A2(n_152), .B1(n_345), .B2(n_497), .C(n_872), .Y(n_916) );
INVx1_ASAP7_75t_L g1303 ( .A(n_17), .Y(n_1303) );
INVxp33_ASAP7_75t_L g831 ( .A(n_18), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_18), .A2(n_133), .B1(n_587), .B2(n_588), .C(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_19), .A2(n_97), .B1(n_491), .B2(n_1041), .Y(n_1040) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_19), .Y(n_1065) );
INVx1_ASAP7_75t_L g1044 ( .A(n_20), .Y(n_1044) );
AO221x2_ASAP7_75t_L g1245 ( .A1(n_21), .A2(n_176), .B1(n_1125), .B2(n_1246), .C(n_1248), .Y(n_1245) );
INVxp33_ASAP7_75t_L g909 ( .A(n_22), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_22), .A2(n_92), .B1(n_920), .B2(n_921), .Y(n_919) );
INVx2_ASAP7_75t_L g292 ( .A(n_23), .Y(n_292) );
OR2x2_ASAP7_75t_L g306 ( .A(n_23), .B(n_290), .Y(n_306) );
INVx1_ASAP7_75t_L g878 ( .A(n_24), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_25), .A2(n_98), .B1(n_314), .B2(n_1297), .Y(n_1296) );
OAI221xp5_ASAP7_75t_L g1327 ( .A1(n_25), .A2(n_98), .B1(n_624), .B2(n_625), .C(n_834), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_26), .A2(n_43), .B1(n_501), .B2(n_774), .C(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g815 ( .A(n_26), .Y(n_815) );
INVx1_ASAP7_75t_L g941 ( .A(n_27), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_28), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_29), .A2(n_129), .B1(n_490), .B2(n_671), .Y(n_1034) );
INVxp33_ASAP7_75t_SL g1054 ( .A(n_29), .Y(n_1054) );
OR2x2_ASAP7_75t_L g282 ( .A(n_30), .B(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g286 ( .A(n_30), .Y(n_286) );
BUFx2_ASAP7_75t_L g374 ( .A(n_30), .Y(n_374) );
INVx1_ASAP7_75t_L g386 ( .A(n_30), .Y(n_386) );
INVxp33_ASAP7_75t_L g908 ( .A(n_31), .Y(n_908) );
AOI21xp33_ASAP7_75t_L g925 ( .A1(n_31), .A2(n_487), .B(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g1042 ( .A(n_32), .Y(n_1042) );
INVx1_ASAP7_75t_L g1312 ( .A(n_33), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_34), .A2(n_143), .B1(n_554), .B2(n_555), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_34), .A2(n_130), .B1(n_515), .B2(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g895 ( .A(n_35), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_36), .A2(n_108), .B1(n_495), .B2(n_496), .C(n_497), .Y(n_494) );
INVx1_ASAP7_75t_L g539 ( .A(n_36), .Y(n_539) );
INVxp33_ASAP7_75t_L g1387 ( .A(n_37), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_37), .A2(n_150), .B1(n_1412), .B2(n_1413), .Y(n_1411) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_38), .Y(n_467) );
OAI221xp5_ASAP7_75t_SL g308 ( .A1(n_39), .A2(n_218), .B1(n_309), .B2(n_314), .C(n_318), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_39), .A2(n_218), .B1(n_407), .B2(n_414), .C(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g850 ( .A(n_40), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_41), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_42), .A2(n_139), .B1(n_343), .B2(n_346), .C(n_350), .Y(n_342) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_42), .Y(n_437) );
INVx1_ASAP7_75t_L g819 ( .A(n_43), .Y(n_819) );
INVx1_ASAP7_75t_L g797 ( .A(n_44), .Y(n_797) );
INVx1_ASAP7_75t_L g1128 ( .A(n_45), .Y(n_1128) );
INVx1_ASAP7_75t_L g1045 ( .A(n_46), .Y(n_1045) );
INVx1_ASAP7_75t_L g729 ( .A(n_47), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_48), .A2(n_189), .B1(n_791), .B2(n_793), .Y(n_1310) );
INVxp67_ASAP7_75t_SL g1318 ( .A(n_48), .Y(n_1318) );
AOI221xp5_ASAP7_75t_SL g484 ( .A1(n_49), .A2(n_64), .B1(n_333), .B2(n_485), .C(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g517 ( .A(n_49), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_50), .A2(n_88), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_50), .A2(n_183), .B1(n_671), .B2(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g481 ( .A(n_51), .Y(n_481) );
INVx1_ASAP7_75t_L g1308 ( .A(n_52), .Y(n_1308) );
INVx1_ASAP7_75t_L g479 ( .A(n_53), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_54), .Y(n_642) );
INVx1_ASAP7_75t_L g341 ( .A(n_55), .Y(n_341) );
INVxp33_ASAP7_75t_L g906 ( .A(n_56), .Y(n_906) );
NAND2xp33_ASAP7_75t_SL g923 ( .A(n_56), .B(n_924), .Y(n_923) );
INVxp33_ASAP7_75t_L g1363 ( .A(n_57), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_57), .A2(n_82), .B1(n_753), .B2(n_1018), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_58), .A2(n_216), .B1(n_491), .B2(n_1299), .C(n_1301), .Y(n_1298) );
INVxp33_ASAP7_75t_L g1333 ( .A(n_58), .Y(n_1333) );
INVx1_ASAP7_75t_L g1292 ( .A(n_59), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_60), .A2(n_193), .B1(n_618), .B2(n_619), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_60), .Y(n_683) );
INVx1_ASAP7_75t_L g1129 ( .A(n_61), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_62), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_63), .A2(n_205), .B1(n_713), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g745 ( .A(n_63), .Y(n_745) );
INVx1_ASAP7_75t_L g514 ( .A(n_64), .Y(n_514) );
INVx1_ASAP7_75t_L g931 ( .A(n_65), .Y(n_931) );
INVxp67_ASAP7_75t_L g996 ( .A(n_66), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_66), .A2(n_170), .B1(n_496), .B2(n_497), .C(n_872), .Y(n_1024) );
XOR2x2_ASAP7_75t_L g549 ( .A(n_67), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g708 ( .A(n_68), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_68), .A2(n_93), .B1(n_490), .B2(n_735), .C(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g1354 ( .A(n_69), .Y(n_1354) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_70), .A2(n_210), .B1(n_472), .B2(n_474), .C(n_477), .Y(n_471) );
INVx1_ASAP7_75t_L g528 ( .A(n_70), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_71), .Y(n_707) );
AO221x1_ASAP7_75t_L g1106 ( .A1(n_72), .A2(n_111), .B1(n_1095), .B2(n_1099), .C(n_1107), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_73), .A2(n_135), .B1(n_281), .B2(n_621), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_73), .Y(n_681) );
INVx1_ASAP7_75t_L g1251 ( .A(n_74), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_74), .A2(n_1338), .B1(n_1341), .B2(n_1434), .Y(n_1337) );
AO22x2_ASAP7_75t_L g1341 ( .A1(n_74), .A2(n_1251), .B1(n_1342), .B2(n_1433), .Y(n_1341) );
INVxp67_ASAP7_75t_L g1003 ( .A(n_75), .Y(n_1003) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_76), .A2(n_164), .B1(n_625), .B2(n_834), .C(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g927 ( .A(n_76), .Y(n_927) );
INVx1_ASAP7_75t_L g367 ( .A(n_77), .Y(n_367) );
AO221x1_ASAP7_75t_L g1113 ( .A1(n_78), .A2(n_159), .B1(n_1095), .B2(n_1099), .C(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1116 ( .A(n_79), .Y(n_1116) );
INVx1_ASAP7_75t_L g290 ( .A(n_80), .Y(n_290) );
INVx1_ASAP7_75t_L g335 ( .A(n_80), .Y(n_335) );
INVx1_ASAP7_75t_L g1070 ( .A(n_81), .Y(n_1070) );
INVx1_ASAP7_75t_L g1353 ( .A(n_82), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_83), .A2(n_245), .B1(n_732), .B2(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g801 ( .A(n_83), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_84), .A2(n_112), .B1(n_834), .B2(n_835), .C(n_901), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_84), .A2(n_112), .B1(n_772), .B2(n_961), .Y(n_1022) );
INVx1_ASAP7_75t_L g478 ( .A(n_85), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_85), .A2(n_210), .B1(n_523), .B2(n_525), .C(n_527), .Y(n_522) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_86), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_86), .A2(n_200), .B1(n_345), .B2(n_495), .C(n_497), .Y(n_865) );
INVx1_ASAP7_75t_L g976 ( .A(n_87), .Y(n_976) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_88), .A2(n_157), .B1(n_485), .B2(n_497), .C(n_968), .Y(n_967) );
INVxp33_ASAP7_75t_SL g828 ( .A(n_89), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_89), .A2(n_107), .B1(n_496), .B2(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_90), .A2(n_227), .B1(n_949), .B2(n_954), .Y(n_953) );
INVxp67_ASAP7_75t_L g966 ( .A(n_90), .Y(n_966) );
INVxp33_ASAP7_75t_SL g943 ( .A(n_91), .Y(n_943) );
AOI21xp33_ASAP7_75t_L g964 ( .A1(n_91), .A2(n_741), .B(n_869), .Y(n_964) );
INVxp33_ASAP7_75t_L g904 ( .A(n_92), .Y(n_904) );
INVx1_ASAP7_75t_L g703 ( .A(n_93), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_94), .A2(n_214), .B1(n_1095), .B2(n_1099), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_95), .A2(n_590), .B(n_592), .C(n_594), .Y(n_589) );
INVx1_ASAP7_75t_L g504 ( .A(n_96), .Y(n_504) );
INVxp33_ASAP7_75t_L g1058 ( .A(n_97), .Y(n_1058) );
INVx1_ASAP7_75t_L g1035 ( .A(n_100), .Y(n_1035) );
INVx1_ASAP7_75t_L g846 ( .A(n_101), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_101), .A2(n_163), .B1(n_671), .B2(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g1111 ( .A(n_102), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_103), .A2(n_154), .B1(n_355), .B2(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g441 ( .A(n_103), .Y(n_441) );
INVx1_ASAP7_75t_L g253 ( .A(n_104), .Y(n_253) );
INVx1_ASAP7_75t_L g896 ( .A(n_106), .Y(n_896) );
INVxp33_ASAP7_75t_SL g832 ( .A(n_107), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_109), .Y(n_581) );
INVxp67_ASAP7_75t_SL g937 ( .A(n_110), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_110), .A2(n_187), .B1(n_309), .B2(n_961), .C(n_962), .Y(n_960) );
XNOR2x1_ASAP7_75t_L g982 ( .A(n_111), .B(n_983), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_113), .A2(n_197), .B1(n_1083), .B2(n_1091), .Y(n_1082) );
INVx1_ASAP7_75t_L g1108 ( .A(n_114), .Y(n_1108) );
INVx1_ASAP7_75t_L g1006 ( .A(n_115), .Y(n_1006) );
INVx1_ASAP7_75t_L g784 ( .A(n_116), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_116), .A2(n_156), .B1(n_723), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_117), .A2(n_138), .B1(n_717), .B2(n_719), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_117), .A2(n_196), .B1(n_352), .B2(n_575), .C(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_118), .A2(n_206), .B1(n_806), .B2(n_952), .Y(n_951) );
INVxp33_ASAP7_75t_L g975 ( .A(n_118), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_119), .A2(n_179), .B1(n_1095), .B2(n_1099), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_120), .A2(n_247), .B1(n_1083), .B2(n_1091), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_121), .A2(n_228), .B1(n_791), .B2(n_793), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_121), .A2(n_131), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g821 ( .A(n_122), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_123), .A2(n_213), .B1(n_407), .B2(n_624), .C(n_625), .Y(n_623) );
OAI222xp33_ASAP7_75t_L g662 ( .A1(n_123), .A2(n_135), .B1(n_213), .B2(n_503), .C1(n_663), .C2(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g898 ( .A(n_124), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_125), .A2(n_180), .B1(n_314), .B2(n_772), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_125), .A2(n_180), .B1(n_625), .B2(n_834), .C(n_901), .Y(n_1055) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_126), .A2(n_575), .B(n_577), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_127), .A2(n_196), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_127), .A2(n_138), .B1(n_752), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g1249 ( .A(n_128), .Y(n_1249) );
INVxp33_ASAP7_75t_L g1050 ( .A(n_129), .Y(n_1050) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_130), .A2(n_145), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_131), .A2(n_140), .B1(n_352), .B2(n_786), .C(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g1365 ( .A(n_132), .Y(n_1365) );
INVxp33_ASAP7_75t_L g829 ( .A(n_133), .Y(n_829) );
INVxp33_ASAP7_75t_L g1348 ( .A(n_134), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_134), .A2(n_148), .B1(n_677), .B2(n_735), .Y(n_1431) );
INVx1_ASAP7_75t_L g1012 ( .A(n_136), .Y(n_1012) );
INVx1_ASAP7_75t_L g1358 ( .A(n_137), .Y(n_1358) );
INVx1_ASAP7_75t_L g432 ( .A(n_139), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_140), .A2(n_228), .B1(n_515), .B2(n_804), .Y(n_803) );
INVxp33_ASAP7_75t_SL g944 ( .A(n_141), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_141), .A2(n_199), .B1(n_328), .B2(n_677), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_142), .A2(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g595 ( .A(n_142), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_143), .A2(n_145), .B1(n_381), .B2(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g796 ( .A(n_144), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_144), .A2(n_175), .B1(n_806), .B2(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g1046 ( .A(n_146), .Y(n_1046) );
INVxp33_ASAP7_75t_L g1345 ( .A(n_148), .Y(n_1345) );
OAI221xp5_ASAP7_75t_L g833 ( .A1(n_149), .A2(n_246), .B1(n_414), .B2(n_834), .C(n_835), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_149), .A2(n_246), .B1(n_309), .B2(n_876), .Y(n_875) );
INVxp33_ASAP7_75t_L g1393 ( .A(n_150), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_151), .A2(n_219), .B1(n_1406), .B2(n_1408), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_151), .A2(n_219), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
INVxp33_ASAP7_75t_L g892 ( .A(n_152), .Y(n_892) );
INVx1_ASAP7_75t_L g319 ( .A(n_153), .Y(n_319) );
INVx1_ASAP7_75t_L g426 ( .A(n_154), .Y(n_426) );
INVx1_ASAP7_75t_L g726 ( .A(n_155), .Y(n_726) );
INVx1_ASAP7_75t_L g795 ( .A(n_156), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_157), .A2(n_183), .B1(n_439), .B2(n_806), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_158), .A2(n_235), .B1(n_495), .B2(n_496), .C(n_497), .Y(n_1309) );
INVxp33_ASAP7_75t_SL g1321 ( .A(n_158), .Y(n_1321) );
INVx1_ASAP7_75t_L g823 ( .A(n_159), .Y(n_823) );
INVx1_ASAP7_75t_L g1295 ( .A(n_160), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_161), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_161), .B(n_253), .Y(n_1090) );
AND3x2_ASAP7_75t_L g1098 ( .A(n_161), .B(n_253), .C(n_1087), .Y(n_1098) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_162), .Y(n_569) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_163), .Y(n_841) );
INVx1_ASAP7_75t_L g928 ( .A(n_164), .Y(n_928) );
INVxp33_ASAP7_75t_L g1395 ( .A(n_165), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_165), .A2(n_178), .B1(n_1408), .B2(n_1416), .Y(n_1415) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_166), .A2(n_204), .B1(n_558), .B2(n_564), .C(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g593 ( .A(n_166), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_167), .Y(n_637) );
INVx2_ASAP7_75t_L g266 ( .A(n_168), .Y(n_266) );
INVx1_ASAP7_75t_L g482 ( .A(n_169), .Y(n_482) );
INVxp33_ASAP7_75t_L g1004 ( .A(n_170), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_171), .A2(n_221), .B1(n_333), .B2(n_652), .C(n_1018), .Y(n_1033) );
INVxp33_ASAP7_75t_L g1051 ( .A(n_171), .Y(n_1051) );
INVx1_ASAP7_75t_L g608 ( .A(n_172), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_173), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_174), .Y(n_644) );
INVx1_ASAP7_75t_L g770 ( .A(n_175), .Y(n_770) );
INVx1_ASAP7_75t_L g1304 ( .A(n_177), .Y(n_1304) );
INVx1_ASAP7_75t_L g1375 ( .A(n_178), .Y(n_1375) );
INVx1_ASAP7_75t_L g1007 ( .A(n_181), .Y(n_1007) );
INVx1_ASAP7_75t_L g1087 ( .A(n_182), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_184), .A2(n_238), .B1(n_302), .B2(n_497), .C(n_1039), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_184), .Y(n_1063) );
INVx1_ASAP7_75t_L g700 ( .A(n_185), .Y(n_700) );
XNOR2x1_ASAP7_75t_L g933 ( .A(n_186), .B(n_934), .Y(n_933) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_187), .Y(n_938) );
AOI22x1_ASAP7_75t_L g882 ( .A1(n_188), .A2(n_883), .B1(n_884), .B2(n_932), .Y(n_882) );
INVx1_ASAP7_75t_L g932 ( .A(n_188), .Y(n_932) );
INVxp33_ASAP7_75t_L g1320 ( .A(n_189), .Y(n_1320) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_190), .Y(n_628) );
INVx1_ASAP7_75t_L g1313 ( .A(n_191), .Y(n_1313) );
INVx1_ASAP7_75t_L g853 ( .A(n_192), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_193), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_194), .Y(n_645) );
INVx1_ASAP7_75t_L g268 ( .A(n_195), .Y(n_268) );
INVx2_ASAP7_75t_L g388 ( .A(n_195), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g1103 ( .A1(n_198), .A2(n_215), .B1(n_1083), .B2(n_1091), .Y(n_1103) );
INVxp33_ASAP7_75t_SL g940 ( .A(n_199), .Y(n_940) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_200), .Y(n_845) );
INVx1_ASAP7_75t_L g1115 ( .A(n_201), .Y(n_1115) );
XOR2xp5_ASAP7_75t_L g1288 ( .A(n_202), .B(n_1289), .Y(n_1288) );
XOR2x1_ASAP7_75t_L g693 ( .A(n_203), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g613 ( .A(n_204), .Y(n_613) );
INVx1_ASAP7_75t_L g758 ( .A(n_205), .Y(n_758) );
INVxp67_ASAP7_75t_L g959 ( .A(n_206), .Y(n_959) );
INVxp33_ASAP7_75t_L g990 ( .A(n_207), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_207), .A2(n_208), .B1(n_333), .B2(n_487), .C(n_1018), .Y(n_1017) );
INVxp33_ASAP7_75t_L g988 ( .A(n_208), .Y(n_988) );
INVxp33_ASAP7_75t_L g891 ( .A(n_209), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_211), .A2(n_225), .B1(n_490), .B2(n_491), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_211), .A2(n_225), .B1(n_511), .B2(n_512), .C(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g851 ( .A(n_212), .Y(n_851) );
INVxp33_ASAP7_75t_L g1330 ( .A(n_216), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_217), .Y(n_634) );
INVx1_ASAP7_75t_L g1011 ( .A(n_220), .Y(n_1011) );
INVxp33_ASAP7_75t_L g1053 ( .A(n_221), .Y(n_1053) );
INVx1_ASAP7_75t_L g1088 ( .A(n_222), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_222), .B(n_1086), .Y(n_1093) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_223), .A2(n_331), .B(n_333), .Y(n_330) );
INVxp33_ASAP7_75t_L g394 ( .A(n_223), .Y(n_394) );
INVxp33_ASAP7_75t_L g399 ( .A(n_224), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_226), .Y(n_1014) );
INVxp33_ASAP7_75t_L g974 ( .A(n_227), .Y(n_974) );
AO22x1_ASAP7_75t_L g1133 ( .A1(n_229), .A2(n_234), .B1(n_1099), .B2(n_1134), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_230), .A2(n_331), .B(n_741), .Y(n_780) );
INVx1_ASAP7_75t_L g818 ( .A(n_230), .Y(n_818) );
INVx1_ASAP7_75t_L g899 ( .A(n_231), .Y(n_899) );
INVx2_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AO22x1_ASAP7_75t_L g1135 ( .A1(n_233), .A2(n_237), .B1(n_1083), .B2(n_1091), .Y(n_1135) );
INVxp67_ASAP7_75t_L g1317 ( .A(n_235), .Y(n_1317) );
INVx1_ASAP7_75t_L g363 ( .A(n_236), .Y(n_363) );
INVxp33_ASAP7_75t_SL g1060 ( .A(n_238), .Y(n_1060) );
INVx1_ASAP7_75t_L g854 ( .A(n_239), .Y(n_854) );
BUFx3_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
INVx1_ASAP7_75t_L g324 ( .A(n_240), .Y(n_324) );
BUFx3_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
INVx1_ASAP7_75t_L g304 ( .A(n_241), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_242), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_243), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_244), .Y(n_779) );
INVx1_ASAP7_75t_L g800 ( .A(n_245), .Y(n_800) );
INVxp33_ASAP7_75t_L g987 ( .A(n_248), .Y(n_987) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_1074), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_251), .B(n_257), .Y(n_1340) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_SL g1336 ( .A(n_252), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_252), .B(n_254), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_254), .B(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x6_ASAP7_75t_L g1372 ( .A(n_259), .B(n_286), .Y(n_1372) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g531 ( .A(n_260), .B(n_268), .Y(n_531) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g421 ( .A(n_261), .B(n_422), .Y(n_421) );
INVx8_ASAP7_75t_L g1364 ( .A(n_262), .Y(n_1364) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_267), .Y(n_262) );
OR2x2_ASAP7_75t_L g281 ( .A(n_263), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g425 ( .A(n_263), .Y(n_425) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_263), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_263), .A2(n_569), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_263), .Y(n_1002) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_263), .Y(n_1010) );
OR2x6_ASAP7_75t_L g1367 ( .A(n_263), .B(n_1347), .Y(n_1367) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x4_ASAP7_75t_L g383 ( .A(n_265), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g392 ( .A(n_265), .Y(n_392) );
AND2x2_ASAP7_75t_L g398 ( .A(n_265), .B(n_266), .Y(n_398) );
INVx2_ASAP7_75t_L g403 ( .A(n_265), .Y(n_403) );
INVx1_ASAP7_75t_L g431 ( .A(n_265), .Y(n_431) );
INVx2_ASAP7_75t_L g384 ( .A(n_266), .Y(n_384) );
INVx1_ASAP7_75t_L g405 ( .A(n_266), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_266), .Y(n_412) );
INVx1_ASAP7_75t_L g430 ( .A(n_266), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_266), .B(n_403), .Y(n_436) );
AND2x4_ASAP7_75t_L g1357 ( .A(n_267), .B(n_412), .Y(n_1357) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B1(n_761), .B2(n_762), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B1(n_692), .B2(n_760), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
XNOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_463), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
XNOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_462), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_375), .Y(n_277) );
AOI21xp33_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_298), .B(n_299), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_279), .A2(n_372), .B1(n_768), .B2(n_797), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_279), .A2(n_911), .B1(n_912), .B2(n_931), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_279), .A2(n_911), .B1(n_957), .B2(n_976), .Y(n_956) );
AOI21xp33_ASAP7_75t_SL g1013 ( .A1(n_279), .A2(n_1014), .B(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_279), .A2(n_911), .B1(n_1031), .B2(n_1046), .Y(n_1030) );
AOI21xp33_ASAP7_75t_L g1291 ( .A1(n_279), .A2(n_1292), .B(n_1293), .Y(n_1291) );
INVx5_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g725 ( .A(n_280), .Y(n_725) );
INVx1_ASAP7_75t_L g879 ( .A(n_280), .Y(n_879) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx2_ASAP7_75t_L g540 ( .A(n_281), .Y(n_540) );
INVx3_ASAP7_75t_L g413 ( .A(n_282), .Y(n_413) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x4_ASAP7_75t_L g1432 ( .A(n_286), .B(n_334), .Y(n_1432) );
INVx2_ASAP7_75t_L g503 ( .A(n_287), .Y(n_503) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_293), .Y(n_287) );
AND2x4_ASAP7_75t_L g310 ( .A(n_288), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_288), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g360 ( .A(n_288), .Y(n_360) );
AND2x4_ASAP7_75t_L g480 ( .A(n_288), .B(n_311), .Y(n_480) );
BUFx2_ASAP7_75t_L g567 ( .A(n_288), .Y(n_567) );
AND2x2_ASAP7_75t_L g733 ( .A(n_288), .B(n_316), .Y(n_733) );
AND2x4_ASAP7_75t_L g877 ( .A(n_288), .B(n_316), .Y(n_877) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g334 ( .A(n_291), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g353 ( .A(n_292), .B(n_335), .Y(n_353) );
INVx1_ASAP7_75t_L g1377 ( .A(n_292), .Y(n_1377) );
HB1xp67_ASAP7_75t_L g1380 ( .A(n_292), .Y(n_1380) );
INVx1_ASAP7_75t_L g1386 ( .A(n_292), .Y(n_1386) );
INVx6_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
BUFx2_ASAP7_75t_L g587 ( .A(n_293), .Y(n_587) );
INVx2_ASAP7_75t_L g754 ( .A(n_293), .Y(n_754) );
AND2x4_ASAP7_75t_L g1388 ( .A(n_293), .B(n_1379), .Y(n_1388) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g317 ( .A(n_294), .Y(n_317) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g340 ( .A(n_295), .B(n_297), .Y(n_340) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g329 ( .A(n_297), .B(n_324), .Y(n_329) );
AOI31xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_336), .A3(n_362), .B(n_371), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B(n_308), .Y(n_300) );
AOI211xp5_ASAP7_75t_L g728 ( .A1(n_301), .A2(n_729), .B(n_730), .C(n_734), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_301), .A2(n_364), .B1(n_795), .B2(n_796), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_301), .A2(n_364), .B1(n_895), .B2(n_898), .Y(n_929) );
AOI21xp33_ASAP7_75t_L g958 ( .A1(n_301), .A2(n_959), .B(n_960), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_301), .A2(n_1006), .B1(n_1017), .B2(n_1019), .C(n_1022), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1032 ( .A1(n_301), .A2(n_1033), .B1(n_1034), .B2(n_1035), .C(n_1036), .Y(n_1032) );
AOI211xp5_ASAP7_75t_L g1294 ( .A1(n_301), .A2(n_1295), .B(n_1296), .C(n_1298), .Y(n_1294) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
BUFx3_ASAP7_75t_L g490 ( .A(n_302), .Y(n_490) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_302), .Y(n_1021) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
BUFx2_ASAP7_75t_L g496 ( .A(n_303), .Y(n_496) );
INVx2_ASAP7_75t_SL g576 ( .A(n_303), .Y(n_576) );
BUFx3_ASAP7_75t_L g585 ( .A(n_303), .Y(n_585) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_303), .Y(n_677) );
AND2x6_ASAP7_75t_L g1394 ( .A(n_303), .B(n_1391), .Y(n_1394) );
INVx1_ASAP7_75t_L g325 ( .A(n_304), .Y(n_325) );
AND2x4_ASAP7_75t_L g338 ( .A(n_305), .B(n_339), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_305), .A2(n_315), .B1(n_471), .B2(n_480), .C1(n_481), .C2(n_482), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_305), .A2(n_553), .B(n_556), .Y(n_552) );
AND2x2_ASAP7_75t_L g863 ( .A(n_305), .B(n_345), .Y(n_863) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g365 ( .A(n_306), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g369 ( .A(n_306), .B(n_370), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_SL g650 ( .A1(n_306), .A2(n_651), .B(n_656), .C(n_661), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_307), .A2(n_367), .B1(n_443), .B2(n_446), .Y(n_442) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g564 ( .A(n_311), .Y(n_564) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g1382 ( .A(n_313), .Y(n_1382) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g565 ( .A(n_316), .Y(n_565) );
INVx2_ASAP7_75t_L g665 ( .A(n_316), .Y(n_665) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x6_ASAP7_75t_L g1376 ( .A(n_317), .B(n_1377), .Y(n_1376) );
OAI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_326), .C(n_330), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_319), .A2(n_378), .B1(n_379), .B2(n_389), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g962 ( .A1(n_320), .A2(n_941), .B(n_963), .C(n_964), .Y(n_962) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g558 ( .A(n_321), .Y(n_558) );
INVx1_ASAP7_75t_L g737 ( .A(n_321), .Y(n_737) );
BUFx4f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g571 ( .A(n_322), .Y(n_571) );
INVx1_ASAP7_75t_L g674 ( .A(n_322), .Y(n_674) );
BUFx2_ASAP7_75t_L g778 ( .A(n_322), .Y(n_778) );
INVx1_ASAP7_75t_L g1302 ( .A(n_322), .Y(n_1302) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
OR2x2_ASAP7_75t_L g366 ( .A(n_323), .B(n_325), .Y(n_366) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g775 ( .A(n_327), .Y(n_775) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_328), .Y(n_671) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
INVx2_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
INVx1_ASAP7_75t_L g492 ( .A(n_329), .Y(n_492) );
INVx1_ASAP7_75t_L g655 ( .A(n_329), .Y(n_655) );
BUFx3_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g488 ( .A(n_332), .Y(n_488) );
INVx1_ASAP7_75t_L g500 ( .A(n_332), .Y(n_500) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_332), .Y(n_562) );
INVx1_ASAP7_75t_L g573 ( .A(n_332), .Y(n_573) );
INVx2_ASAP7_75t_SL g869 ( .A(n_332), .Y(n_869) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_332), .Y(n_971) );
INVx2_ASAP7_75t_L g1397 ( .A(n_332), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g588 ( .A(n_334), .Y(n_588) );
INVx2_ASAP7_75t_L g741 ( .A(n_334), .Y(n_741) );
INVx2_ASAP7_75t_SL g1306 ( .A(n_334), .Y(n_1306) );
INVx1_ASAP7_75t_L g1399 ( .A(n_335), .Y(n_1399) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B1(n_342), .B2(n_354), .C(n_358), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_337), .A2(n_358), .B1(n_1012), .B2(n_1024), .C(n_1025), .Y(n_1023) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g744 ( .A(n_338), .Y(n_744) );
INVx2_ASAP7_75t_SL g783 ( .A(n_338), .Y(n_783) );
INVx1_ASAP7_75t_L g915 ( .A(n_338), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_338), .A2(n_358), .B1(n_1038), .B2(n_1040), .C(n_1042), .Y(n_1037) );
INVx2_ASAP7_75t_SL g486 ( .A(n_339), .Y(n_486) );
BUFx3_ASAP7_75t_L g495 ( .A(n_339), .Y(n_495) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_339), .Y(n_660) );
AND2x4_ASAP7_75t_L g972 ( .A(n_339), .B(n_567), .Y(n_972) );
BUFx4f_ASAP7_75t_L g1018 ( .A(n_339), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_340), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_341), .A2(n_363), .B1(n_450), .B2(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_345), .A2(n_361), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g555 ( .A(n_345), .Y(n_555) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_349), .Y(n_361) );
INVx2_ASAP7_75t_L g750 ( .A(n_349), .Y(n_750) );
AND2x4_ASAP7_75t_L g1389 ( .A(n_349), .B(n_1390), .Y(n_1389) );
BUFx6f_ASAP7_75t_L g1422 ( .A(n_349), .Y(n_1422) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
BUFx3_ASAP7_75t_L g498 ( .A(n_353), .Y(n_498) );
INVx2_ASAP7_75t_L g579 ( .A(n_353), .Y(n_579) );
INVx1_ASAP7_75t_L g1428 ( .A(n_353), .Y(n_1428) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g557 ( .A(n_357), .Y(n_557) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_357), .Y(n_735) );
INVx1_ASAP7_75t_L g922 ( .A(n_357), .Y(n_922) );
AND2x6_ASAP7_75t_L g1384 ( .A(n_357), .B(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1425 ( .A(n_357), .Y(n_1425) );
AOI21xp33_ASAP7_75t_L g483 ( .A1(n_358), .A2(n_484), .B(n_489), .Y(n_483) );
INVx1_ASAP7_75t_L g661 ( .A(n_358), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_358), .A2(n_743), .B1(n_745), .B2(n_746), .C(n_751), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_358), .A2(n_782), .B1(n_784), .B2(n_785), .C(n_790), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_358), .A2(n_782), .B1(n_854), .B2(n_865), .C(n_866), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_358), .A2(n_896), .B1(n_914), .B2(n_916), .C(n_917), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_358), .A2(n_914), .B1(n_1308), .B2(n_1309), .C(n_1310), .Y(n_1307) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g664 ( .A(n_360), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g789 ( .A(n_361), .Y(n_789) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_361), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_367), .B2(n_368), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_364), .A2(n_368), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_364), .A2(n_850), .B1(n_853), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_364), .A2(n_368), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_364), .A2(n_368), .B1(n_1007), .B2(n_1011), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_364), .A2(n_368), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g1311 ( .A1(n_364), .A2(n_368), .B1(n_1312), .B2(n_1313), .Y(n_1311) );
INVx6_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g473 ( .A(n_366), .Y(n_473) );
INVx1_ASAP7_75t_L g739 ( .A(n_366), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_368), .A2(n_770), .B(n_771), .C(n_773), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_368), .A2(n_851), .B1(n_871), .B2(n_873), .C(n_875), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_368), .B(n_899), .Y(n_930) );
INVx4_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g476 ( .A(n_370), .Y(n_476) );
INVx1_ASAP7_75t_L g874 ( .A(n_370), .Y(n_874) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g858 ( .A(n_373), .Y(n_858) );
AND2x4_ASAP7_75t_L g1398 ( .A(n_373), .B(n_1399), .Y(n_1398) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x6_ASAP7_75t_L g420 ( .A(n_374), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g507 ( .A(n_374), .Y(n_507) );
NOR3xp33_ASAP7_75t_SL g375 ( .A(n_376), .B(n_406), .C(n_419), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_393), .Y(n_376) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g704 ( .A(n_380), .Y(n_704) );
BUFx2_ASAP7_75t_L g816 ( .A(n_380), .Y(n_816) );
BUFx2_ASAP7_75t_L g905 ( .A(n_380), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_380), .A2(n_389), .B1(n_987), .B2(n_988), .Y(n_986) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_380), .Y(n_1331) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_385), .Y(n_380) );
BUFx3_ASAP7_75t_L g807 ( .A(n_381), .Y(n_807) );
INVx1_ASAP7_75t_L g1325 ( .A(n_381), .Y(n_1325) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
BUFx6f_ASAP7_75t_L g1404 ( .A(n_382), .Y(n_1404) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
INVx1_ASAP7_75t_L g1351 ( .A(n_383), .Y(n_1351) );
INVx1_ASAP7_75t_L g1414 ( .A(n_383), .Y(n_1414) );
AND2x4_ASAP7_75t_L g391 ( .A(n_384), .B(n_392), .Y(n_391) );
AND2x6_ASAP7_75t_L g389 ( .A(n_385), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g395 ( .A(n_385), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_385), .B(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_385), .A2(n_510), .B1(n_521), .B2(n_522), .Y(n_509) );
AND2x2_ASAP7_75t_L g591 ( .A(n_385), .B(n_401), .Y(n_591) );
AND2x2_ASAP7_75t_L g596 ( .A(n_385), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g599 ( .A(n_385), .B(n_448), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_385), .B(n_605), .Y(n_611) );
AND2x2_ASAP7_75t_L g820 ( .A(n_385), .B(n_401), .Y(n_820) );
AND2x2_ASAP7_75t_L g992 ( .A(n_385), .B(n_401), .Y(n_992) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g458 ( .A(n_386), .Y(n_458) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
INVx1_ASAP7_75t_L g460 ( .A(n_388), .Y(n_460) );
INVx1_ASAP7_75t_SL g619 ( .A(n_389), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_389), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_389), .A2(n_779), .B1(n_815), .B2(n_816), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_389), .A2(n_816), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_389), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_389), .A2(n_905), .B1(n_940), .B2(n_941), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_389), .A2(n_816), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_389), .A2(n_1303), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_390), .B(n_413), .Y(n_418) );
BUFx2_ASAP7_75t_L g949 ( .A(n_390), .Y(n_949) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_391), .Y(n_520) );
BUFx2_ASAP7_75t_L g548 ( .A(n_391), .Y(n_548) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_391), .Y(n_605) );
INVx1_ASAP7_75t_L g715 ( .A(n_391), .Y(n_715) );
AND2x4_ASAP7_75t_L g1369 ( .A(n_391), .B(n_1370), .Y(n_1369) );
BUFx3_ASAP7_75t_L g1409 ( .A(n_391), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_399), .B2(n_400), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_395), .A2(n_400), .B1(n_707), .B2(n_708), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_395), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_395), .A2(n_820), .B1(n_831), .B2(n_832), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_395), .A2(n_820), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_395), .A2(n_400), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_395), .A2(n_990), .B1(n_991), .B2(n_992), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_395), .A2(n_400), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_395), .A2(n_820), .B1(n_1304), .B2(n_1333), .Y(n_1332) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g597 ( .A(n_397), .Y(n_597) );
INVx2_ASAP7_75t_L g813 ( .A(n_397), .Y(n_813) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_398), .Y(n_516) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g524 ( .A(n_402), .Y(n_524) );
INVx1_ASAP7_75t_L g534 ( .A(n_402), .Y(n_534) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_402), .Y(n_603) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_402), .Y(n_718) );
BUFx2_ASAP7_75t_L g806 ( .A(n_402), .Y(n_806) );
AND2x4_ASAP7_75t_L g1346 ( .A(n_402), .B(n_1347), .Y(n_1346) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g416 ( .A(n_403), .Y(n_416) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g834 ( .A(n_408), .Y(n_834) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2x1_ASAP7_75t_SL g409 ( .A(n_410), .B(n_413), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_412), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_413), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g542 ( .A(n_413), .B(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g544 ( .A(n_413), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g547 ( .A(n_413), .B(n_548), .Y(n_547) );
BUFx4f_ASAP7_75t_L g624 ( .A(n_414), .Y(n_624) );
BUFx4f_ASAP7_75t_L g901 ( .A(n_414), .Y(n_901) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g625 ( .A(n_418), .Y(n_625) );
BUFx2_ASAP7_75t_L g835 ( .A(n_418), .Y(n_835) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .A3(n_433), .B1(n_442), .B2(n_449), .B3(n_455), .Y(n_419) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_420), .Y(n_837) );
OAI33xp33_ASAP7_75t_L g886 ( .A1(n_420), .A2(n_455), .A3(n_887), .B1(n_890), .B2(n_894), .B3(n_897), .Y(n_886) );
OAI33xp33_ASAP7_75t_L g994 ( .A1(n_420), .A2(n_455), .A3(n_995), .B1(n_1000), .B2(n_1005), .B3(n_1008), .Y(n_994) );
OAI33xp33_ASAP7_75t_L g1056 ( .A1(n_420), .A2(n_455), .A3(n_1057), .B1(n_1062), .B2(n_1067), .B3(n_1069), .Y(n_1056) );
OAI33xp33_ASAP7_75t_L g1315 ( .A1(n_420), .A2(n_455), .A3(n_1316), .B1(n_1319), .B2(n_1324), .B3(n_1326), .Y(n_1315) );
INVx1_ASAP7_75t_L g1347 ( .A(n_422), .Y(n_1347) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_432), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g633 ( .A(n_425), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_427), .A2(n_839), .B1(n_895), .B2(n_896), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_427), .A2(n_1042), .B1(n_1044), .B2(n_1059), .Y(n_1069) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g454 ( .A(n_429), .Y(n_454) );
INVx2_ASAP7_75t_L g1061 ( .A(n_429), .Y(n_1061) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_430), .B(n_431), .Y(n_610) );
INVx1_ASAP7_75t_L g546 ( .A(n_431), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_433) );
BUFx2_ASAP7_75t_L g844 ( .A(n_434), .Y(n_844) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g445 ( .A(n_436), .Y(n_445) );
BUFx2_ASAP7_75t_L g640 ( .A(n_436), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_438), .A2(n_443), .B1(n_898), .B2(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g512 ( .A(n_440), .Y(n_512) );
INVx2_ASAP7_75t_SL g536 ( .A(n_440), .Y(n_536) );
INVx4_ASAP7_75t_L g630 ( .A(n_440), .Y(n_630) );
INVx2_ASAP7_75t_SL g720 ( .A(n_440), .Y(n_720) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_440), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_443), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g849 ( .A(n_445), .Y(n_849) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g526 ( .A(n_448), .Y(n_526) );
INVx2_ASAP7_75t_L g641 ( .A(n_448), .Y(n_641) );
INVx2_ASAP7_75t_L g810 ( .A(n_448), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_450), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_452), .A2(n_454), .B1(n_479), .B2(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_452), .A2(n_454), .B1(n_538), .B2(n_539), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g643 ( .A1(n_452), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g840 ( .A(n_452), .Y(n_840) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_452), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_453), .A2(n_839), .B1(n_841), .B2(n_842), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_453), .A2(n_1009), .B1(n_1011), .B2(n_1012), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_453), .A2(n_1009), .B1(n_1308), .B2(n_1312), .Y(n_1326) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g1323 ( .A(n_454), .Y(n_1323) );
OAI33xp33_ASAP7_75t_L g836 ( .A1(n_455), .A2(n_837), .A3(n_838), .B1(n_843), .B2(n_847), .B3(n_852), .Y(n_836) );
CKINVDCx8_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx6_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g1418 ( .A(n_459), .Y(n_1418) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g1361 ( .A(n_460), .Y(n_1361) );
OAI22x1_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_614), .B2(n_691), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
XNOR2x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_549), .Y(n_465) );
XNOR2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_508), .Y(n_468) );
AOI31xp33_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_483), .A3(n_493), .B(n_505), .Y(n_469) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_473), .Y(n_669) );
INVx2_ASAP7_75t_L g684 ( .A(n_473), .Y(n_684) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g756 ( .A(n_476), .Y(n_756) );
INVx2_ASAP7_75t_SL g663 ( .A(n_480), .Y(n_663) );
INVx1_ASAP7_75t_L g731 ( .A(n_480), .Y(n_731) );
INVx2_ASAP7_75t_SL g772 ( .A(n_480), .Y(n_772) );
AOI322xp5_ASAP7_75t_L g918 ( .A1(n_480), .A2(n_733), .A3(n_919), .B1(n_923), .B2(n_925), .C1(n_927), .C2(n_928), .Y(n_918) );
INVx1_ASAP7_75t_L g1297 ( .A(n_480), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_481), .A2(n_482), .B1(n_542), .B2(n_544), .C(n_547), .Y(n_541) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g924 ( .A(n_486), .Y(n_924) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g792 ( .A(n_488), .Y(n_792) );
INVxp67_ASAP7_75t_L g680 ( .A(n_490), .Y(n_680) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g501 ( .A(n_492), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_499), .B1(n_502), .B2(n_504), .Y(n_493) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_498), .A2(n_628), .B1(n_634), .B2(n_673), .C(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_504), .A2(n_530), .B1(n_532), .B2(n_540), .Y(n_529) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_506), .A2(n_551), .B(n_589), .C(n_600), .Y(n_550) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g530 ( .A(n_507), .B(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g688 ( .A(n_507), .Y(n_688) );
AND2x4_ASAP7_75t_L g711 ( .A(n_507), .B(n_531), .Y(n_711) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_507), .B(n_1418), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_507), .B(n_1428), .Y(n_1427) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_529), .C(n_541), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_513) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_515), .Y(n_948) );
INVx1_ASAP7_75t_L g955 ( .A(n_515), .Y(n_955) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g713 ( .A(n_516), .Y(n_713) );
INVx3_ASAP7_75t_L g1407 ( .A(n_516), .Y(n_1407) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g804 ( .A(n_519), .Y(n_804) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AOI322xp5_ASAP7_75t_L g601 ( .A1(n_521), .A2(n_530), .A3(n_581), .B1(n_602), .B2(n_604), .C1(n_606), .C2(n_611), .Y(n_601) );
AOI33xp33_ASAP7_75t_L g709 ( .A1(n_521), .A2(n_710), .A3(n_712), .B1(n_716), .B2(n_721), .B3(n_722), .Y(n_709) );
AOI33xp33_ASAP7_75t_L g802 ( .A1(n_521), .A2(n_530), .A3(n_803), .B1(n_805), .B2(n_808), .B3(n_811), .Y(n_802) );
AOI33xp33_ASAP7_75t_L g945 ( .A1(n_521), .A2(n_946), .A3(n_947), .B1(n_950), .B2(n_951), .B3(n_953), .Y(n_945) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g952 ( .A(n_526), .Y(n_952) );
BUFx2_ASAP7_75t_L g946 ( .A(n_530), .Y(n_946) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g1412 ( .A(n_534), .Y(n_1412) );
INVxp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_540), .A2(n_544), .B1(n_560), .B2(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_542), .A2(n_547), .B(n_613), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_542), .A2(n_697), .B1(n_699), .B2(n_700), .C(n_701), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g799 ( .A1(n_542), .A2(n_544), .B1(n_547), .B2(n_800), .C(n_801), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_542), .A2(n_544), .B1(n_547), .B2(n_937), .C(n_938), .Y(n_936) );
INVx1_ASAP7_75t_L g698 ( .A(n_544), .Y(n_698) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_545), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_547), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g1352 ( .A1(n_548), .A2(n_1353), .B1(n_1354), .B2(n_1355), .C1(n_1358), .C2(n_1359), .Y(n_1352) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_552), .B(n_559), .C(n_568), .D(n_580), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_557), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g793 ( .A(n_557), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_563), .C(n_566), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g652 ( .A(n_562), .Y(n_652) );
INVx1_ASAP7_75t_L g1421 ( .A(n_562), .Y(n_1421) );
BUFx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_572), .C(n_574), .Y(n_568) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g583 ( .A(n_571), .Y(n_583) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g920 ( .A(n_576), .Y(n_920) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_584), .C(n_586), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g658 ( .A(n_585), .Y(n_658) );
INVx1_ASAP7_75t_L g686 ( .A(n_588), .Y(n_686) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g618 ( .A(n_591), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g648 ( .A(n_596), .Y(n_648) );
INVx2_ASAP7_75t_L g621 ( .A(n_599), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_612), .Y(n_600) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_605), .Y(n_723) );
BUFx3_ASAP7_75t_L g635 ( .A(n_609), .Y(n_635) );
INVx2_ASAP7_75t_L g647 ( .A(n_609), .Y(n_647) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g691 ( .A(n_614), .Y(n_691) );
INVx1_ASAP7_75t_L g689 ( .A(n_615), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_622), .C(n_649), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_629), .A2(n_632), .B1(n_668), .B2(n_670), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_630), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_630), .A2(n_848), .B1(n_850), .B2(n_851), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_630), .A2(n_996), .B1(n_997), .B2(n_999), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_641), .B2(n_642), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_637), .A2(n_645), .B1(n_657), .B2(n_659), .Y(n_656) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_641), .A2(n_844), .B1(n_888), .B2(n_889), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_641), .A2(n_997), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_642), .A2(n_644), .B1(n_652), .B2(n_653), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_646), .A2(n_839), .B1(n_853), .B2(n_854), .Y(n_852) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g893 ( .A(n_647), .Y(n_893) );
OAI31xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_662), .A3(n_666), .B(n_687), .Y(n_649) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .B1(n_678), .B2(n_682), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_682) );
BUFx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g787 ( .A(n_677), .Y(n_787) );
INVx2_ASAP7_75t_L g1300 ( .A(n_677), .Y(n_1300) );
CKINVDCx8_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g727 ( .A1(n_688), .A2(n_728), .A3(n_742), .B(n_757), .Y(n_727) );
INVxp67_ASAP7_75t_L g760 ( .A(n_692), .Y(n_760) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_724), .Y(n_694) );
AND4x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_702), .C(n_706), .D(n_709), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_705), .A2(n_707), .B1(n_737), .B2(n_738), .C(n_740), .Y(n_736) );
BUFx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g1401 ( .A(n_711), .B(n_1402), .C(n_1405), .Y(n_1401) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI21xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_727), .Y(n_724) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g1301 ( .A1(n_738), .A2(n_1302), .B1(n_1303), .B2(n_1304), .C(n_1305), .Y(n_1301) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g926 ( .A(n_741), .Y(n_926) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
BUFx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g1041 ( .A(n_754), .Y(n_1041) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_979), .B1(n_980), .B2(n_1073), .Y(n_762) );
INVx1_ASAP7_75t_L g1073 ( .A(n_763), .Y(n_1073) );
XNOR2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_880), .Y(n_763) );
XOR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_822), .Y(n_764) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_821), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_798), .Y(n_766) );
NAND3xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_781), .C(n_794), .Y(n_768) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g968 ( .A(n_775), .Y(n_968) );
OAI21xp5_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_779), .B(n_780), .Y(n_776) );
INVx2_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g1039 ( .A(n_789), .Y(n_1039) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AND4x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .C(n_814), .D(n_817), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_807), .Y(n_1068) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
XNOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_855), .Y(n_824) );
NOR3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_833), .C(n_836), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_830), .Y(n_826) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g998 ( .A(n_849), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_859), .B1(n_878), .B2(n_879), .Y(n_855) );
INVx5_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI31xp33_ASAP7_75t_L g1015 ( .A1(n_857), .A2(n_1016), .A3(n_1023), .B(n_1026), .Y(n_1015) );
AOI31xp33_ASAP7_75t_L g1293 ( .A1(n_857), .A2(n_1294), .A3(n_1307), .B(n_1311), .Y(n_1293) );
BUFx8_ASAP7_75t_SL g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g911 ( .A(n_858), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_864), .C(n_870), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AOI222xp33_ASAP7_75t_L g1374 ( .A1(n_872), .A2(n_1354), .B1(n_1358), .B2(n_1375), .C1(n_1376), .C2(n_1378), .Y(n_1374) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_SL g961 ( .A(n_877), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_933), .B1(n_977), .B2(n_978), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_882), .Y(n_978) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_910), .Y(n_884) );
NOR3xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_900), .C(n_902), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_893), .A2(n_1001), .B1(n_1003), .B2(n_1004), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_907), .Y(n_902) );
NAND4xp25_ASAP7_75t_L g912 ( .A(n_913), .B(n_918), .C(n_929), .D(n_930), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_914), .A2(n_966), .B1(n_967), .B2(n_969), .C(n_972), .Y(n_965) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g977 ( .A(n_933), .Y(n_977) );
AND2x2_ASAP7_75t_L g934 ( .A(n_935), .B(n_956), .Y(n_934) );
AND4x1_ASAP7_75t_L g935 ( .A(n_936), .B(n_939), .C(n_942), .D(n_945), .Y(n_935) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NAND3xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_965), .C(n_973), .Y(n_957) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1027), .B1(n_1071), .B2(n_1072), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
BUFx2_ASAP7_75t_SL g1071 ( .A(n_982), .Y(n_1071) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_1013), .Y(n_983) );
NOR3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_993), .C(n_994), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_997), .A2(n_1068), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_L g1064 ( .A(n_998), .Y(n_1064) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx3_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
BUFx2_ASAP7_75t_SL g1072 ( .A(n_1028), .Y(n_1072) );
XOR2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1070), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1047), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1037), .C(n_1043), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1035), .A2(n_1045), .B1(n_1064), .B2(n_1068), .Y(n_1067) );
NOR3xp33_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1055), .C(n_1056), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1052), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1059), .B1(n_1060), .B2(n_1061), .Y(n_1057) );
OAI22xp33_ASAP7_75t_L g1319 ( .A1(n_1059), .A2(n_1320), .B1(n_1321), .B2(n_1322), .Y(n_1319) );
OAI22xp5_ASAP7_75t_SL g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1064), .A2(n_1295), .B1(n_1313), .B2(n_1325), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1284), .B1(n_1288), .B2(n_1334), .C(n_1337), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1211), .Y(n_1075) );
NOR2xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1193), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1150), .C(n_1179), .Y(n_1077) );
O2A1O1Ixp33_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1117), .B(n_1122), .C(n_1136), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1100), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1080), .B(n_1139), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1080), .B(n_1160), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1080), .B(n_1123), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1080), .B(n_1101), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1080), .B(n_1178), .Y(n_1192) );
OAI332xp33_ASAP7_75t_L g1215 ( .A1(n_1080), .A2(n_1147), .A3(n_1166), .B1(n_1167), .B2(n_1216), .B3(n_1219), .C1(n_1220), .C2(n_1222), .Y(n_1215) );
OAI32xp33_ASAP7_75t_L g1277 ( .A1(n_1080), .A2(n_1208), .A3(n_1233), .B1(n_1263), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1080), .Y(n_1279) );
INVx4_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1081), .B(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1081), .B(n_1139), .Y(n_1147) );
INVx3_ASAP7_75t_L g1165 ( .A(n_1081), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1081), .B(n_1167), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1081), .B(n_1187), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1081), .B(n_1139), .Y(n_1231) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1081), .B(n_1218), .Y(n_1274) );
NAND3xp33_ASAP7_75t_L g1281 ( .A(n_1081), .B(n_1264), .C(n_1275), .Y(n_1281) );
NOR3xp33_ASAP7_75t_L g1282 ( .A(n_1081), .B(n_1161), .C(n_1283), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1094), .Y(n_1081) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1089), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_1085), .B(n_1090), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1088), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_1089), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1090), .B(n_1093), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_1092), .Y(n_1436) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1095), .Y(n_1247) );
AND2x4_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1098), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1096), .B(n_1098), .Y(n_1134) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1097), .B(n_1098), .Y(n_1099) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1099), .Y(n_1126) );
OAI21xp5_ASAP7_75t_L g1144 ( .A1(n_1100), .A2(n_1145), .B(n_1146), .Y(n_1144) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1100), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1100), .B(n_1164), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_1100), .A2(n_1170), .B1(n_1266), .B2(n_1273), .C(n_1274), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1105), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1101), .B(n_1118), .Y(n_1117) );
NOR2x1_ASAP7_75t_L g1160 ( .A(n_1101), .B(n_1161), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1101), .B(n_1161), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1101), .B(n_1186), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1101), .B(n_1156), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1101), .B(n_1225), .Y(n_1224) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1102), .B(n_1105), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1102), .B(n_1120), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1102), .B(n_1155), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1102), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1102), .B(n_1161), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1102), .B(n_1186), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1102), .B(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1105), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1105), .Y(n_1218) );
OAI21xp5_ASAP7_75t_L g1265 ( .A1(n_1105), .A2(n_1221), .B(n_1266), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1113), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1106), .B(n_1121), .Y(n_1120) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1106), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1109), .B1(n_1111), .B2(n_1112), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_1109), .A2(n_1112), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1127 ( .A1(n_1109), .A2(n_1128), .B1(n_1129), .B2(n_1130), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1250 ( .A(n_1109), .Y(n_1250) );
BUFx6f_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1112), .Y(n_1130) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1112), .Y(n_1253) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1113), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1113), .B(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1113), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_1117), .A2(n_1178), .B1(n_1198), .B2(n_1202), .C(n_1203), .Y(n_1197) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1120), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1121), .B(n_1156), .Y(n_1186) );
NAND3xp33_ASAP7_75t_L g1171 ( .A(n_1122), .B(n_1169), .C(n_1172), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1122), .B(n_1170), .Y(n_1240) );
AND2x4_ASAP7_75t_SL g1122 ( .A(n_1123), .B(n_1131), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1123), .B(n_1132), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1123), .B(n_1131), .Y(n_1208) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_1124), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1124), .B(n_1131), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1124), .B(n_1169), .Y(n_1168) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1124), .Y(n_1205) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1131), .B(n_1170), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1131), .B(n_1139), .Y(n_1264) );
CKINVDCx6p67_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1132), .B(n_1139), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1132), .B(n_1188), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_1132), .Y(n_1222) );
OR2x6_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1135), .Y(n_1132) );
O2A1O1Ixp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1142), .B(n_1144), .C(n_1148), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1138), .B(n_1186), .Y(n_1227) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1139), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_1139), .Y(n_1170) );
INVx1_ASAP7_75t_SL g1188 ( .A(n_1139), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
AOI21xp33_ASAP7_75t_SL g1174 ( .A1(n_1142), .A2(n_1175), .B(n_1176), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1142), .B(n_1170), .Y(n_1259) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_1143), .A2(n_1238), .B(n_1239), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1143), .B(n_1214), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1145), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1149), .B(n_1188), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1149), .B(n_1227), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1149), .B(n_1165), .Y(n_1257) );
AOI211xp5_ASAP7_75t_SL g1150 ( .A1(n_1151), .A2(n_1154), .B(n_1157), .C(n_1174), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1152), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g1278 ( .A(n_1153), .B(n_1273), .C(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1155), .B(n_1182), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1155), .B(n_1165), .Y(n_1225) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1155), .Y(n_1242) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1156), .Y(n_1273) );
OAI221xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1162), .B1(n_1163), .B2(n_1168), .C(n_1171), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1161), .B(n_1167), .Y(n_1166) );
AOI222xp33_ASAP7_75t_L g1276 ( .A1(n_1161), .A2(n_1183), .B1(n_1245), .B2(n_1277), .C1(n_1280), .C2(n_1282), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1164), .B(n_1183), .Y(n_1232) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1165), .B(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1165), .B(n_1200), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1165), .B(n_1221), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1167), .B(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1168), .Y(n_1238) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1170), .B(n_1210), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1178), .B(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1178), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1183), .B1(n_1184), .B2(n_1187), .C(n_1189), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1182), .B(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1186), .Y(n_1217) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1187), .Y(n_1271) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_1190), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1191), .Y(n_1233) );
OAI211xp5_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1195), .B(n_1197), .C(n_1206), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_1194), .A2(n_1220), .B1(n_1241), .B2(n_1257), .C(n_1258), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1201), .Y(n_1198) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_1199), .A2(n_1208), .B1(n_1222), .B2(n_1224), .C(n_1226), .Y(n_1223) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1205), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1230 ( .A(n_1205), .B(n_1231), .Y(n_1230) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1205), .Y(n_1235) );
OAI31xp33_ASAP7_75t_L g1260 ( .A1(n_1205), .A2(n_1261), .A3(n_1263), .B(n_1265), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1205), .B(n_1245), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1209), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
AOI21xp5_ASAP7_75t_L g1211 ( .A1(n_1212), .A2(n_1243), .B(n_1254), .Y(n_1211) );
NAND3xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1234), .C(n_1237), .Y(n_1212) );
AOI211xp5_ASAP7_75t_L g1213 ( .A1(n_1214), .A2(n_1215), .B(n_1223), .C(n_1228), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI221xp5_ASAP7_75t_SL g1269 ( .A1(n_1222), .A2(n_1242), .B1(n_1270), .B2(n_1271), .C(n_1272), .Y(n_1269) );
AOI21xp33_ASAP7_75t_SL g1228 ( .A1(n_1229), .A2(n_1232), .B(n_1233), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1231), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
OAI31xp33_ASAP7_75t_L g1255 ( .A1(n_1244), .A2(n_1256), .A3(n_1259), .B(n_1260), .Y(n_1255) );
BUFx3_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1245), .Y(n_1283) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1250), .B1(n_1251), .B2(n_1252), .Y(n_1248) );
HB1xp67_ASAP7_75t_L g1287 ( .A(n_1252), .Y(n_1287) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1267), .C(n_1276), .Y(n_1254) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI21xp33_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .B(n_1275), .Y(n_1267) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_SL g1285 ( .A(n_1286), .Y(n_1285) );
BUFx2_ASAP7_75t_SL g1286 ( .A(n_1287), .Y(n_1286) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1314), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NOR3xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1327), .C(n_1328), .Y(n_1314) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1332), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_1335), .Y(n_1334) );
OAI21xp5_ASAP7_75t_L g1435 ( .A1(n_1336), .A2(n_1436), .B(n_1437), .Y(n_1435) );
BUFx3_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1342), .Y(n_1433) );
AOI221x1_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1371), .B1(n_1373), .B2(n_1398), .C(n_1400), .Y(n_1342) );
NAND4xp25_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1352), .C(n_1362), .D(n_1368), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1346), .B1(n_1348), .B2(n_1349), .Y(n_1344) );
AND2x4_ASAP7_75t_L g1349 ( .A(n_1347), .B(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1361), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1364), .B1(n_1365), .B2(n_1366), .Y(n_1362) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_1365), .A2(n_1384), .B1(n_1387), .B2(n_1388), .C(n_1389), .Y(n_1383) );
INVx5_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
CKINVDCx11_ASAP7_75t_R g1368 ( .A(n_1369), .Y(n_1368) );
CKINVDCx16_ASAP7_75t_R g1371 ( .A(n_1372), .Y(n_1371) );
NAND3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1383), .C(n_1392), .Y(n_1373) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1377), .Y(n_1391) );
AND2x2_ASAP7_75t_SL g1378 ( .A(n_1379), .B(n_1381), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
AND2x4_ASAP7_75t_L g1396 ( .A(n_1385), .B(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_SL g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1392 ( .A1(n_1393), .A2(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1392) );
NAND4xp25_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1410), .C(n_1419), .D(n_1429), .Y(n_1400) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_1407), .Y(n_1416) );
BUFx6f_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
NAND3xp33_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1415), .C(n_1417), .Y(n_1410) );
INVx2_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
NAND3xp33_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1423), .C(n_1426), .Y(n_1419) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx3_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
NAND3xp33_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1431), .C(n_1432), .Y(n_1429) );
HB1xp67_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
endmodule