module fake_jpeg_13685_n_468 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_468);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_468;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_55),
.B(n_65),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_67),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_73),
.Y(n_178)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_33),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_80),
.B(n_83),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_33),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_10),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_102),
.Y(n_168)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_89),
.B(n_8),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_92),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_42),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_31),
.B(n_9),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_31),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_112),
.Y(n_196)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_111),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_19),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_116),
.Y(n_167)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_44),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_118),
.Y(n_183)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_29),
.B1(n_73),
.B2(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_120),
.A2(n_128),
.B1(n_130),
.B2(n_140),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_51),
.B1(n_40),
.B2(n_20),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_51),
.B1(n_40),
.B2(n_48),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_51),
.B1(n_43),
.B2(n_19),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_134),
.A2(n_139),
.B(n_171),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_43),
.B1(n_35),
.B2(n_25),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_62),
.A2(n_53),
.B1(n_48),
.B2(n_46),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_69),
.A2(n_104),
.B1(n_88),
.B2(n_100),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_53),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_143),
.B(n_153),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_57),
.A2(n_52),
.B1(n_47),
.B2(n_20),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_146),
.A2(n_159),
.B1(n_164),
.B2(n_180),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_67),
.B(n_46),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_108),
.A2(n_113),
.B1(n_112),
.B2(n_35),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_52),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_161),
.B(n_186),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_69),
.A2(n_102),
.B1(n_118),
.B2(n_56),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_66),
.A2(n_47),
.B1(n_25),
.B2(n_2),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

AO22x1_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_134),
.B1(n_158),
.B2(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_8),
.C(n_3),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_59),
.A2(n_81),
.B1(n_78),
.B2(n_111),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_176),
.B(n_184),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_3),
.B1(n_7),
.B2(n_71),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_86),
.A2(n_3),
.B1(n_90),
.B2(n_103),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_107),
.B1(n_105),
.B2(n_84),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_181),
.A2(n_182),
.B1(n_137),
.B2(n_127),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_61),
.A2(n_77),
.B1(n_39),
.B2(n_50),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_106),
.A2(n_24),
.B1(n_18),
.B2(n_41),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_107),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_60),
.A2(n_24),
.B1(n_18),
.B2(n_41),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_190),
.B(n_172),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_60),
.A2(n_24),
.B1(n_18),
.B2(n_41),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_107),
.B(n_55),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_107),
.B(n_55),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_197),
.B(n_200),
.Y(n_273)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_160),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_158),
.Y(n_201)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_202),
.B(n_229),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_154),
.C(n_161),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_203),
.B(n_232),
.Y(n_301)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_204),
.Y(n_303)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_123),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_206),
.B(n_209),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_168),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_207),
.B(n_237),
.C(n_248),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_139),
.B(n_136),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_145),
.B(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_210),
.B(n_212),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_150),
.B1(n_156),
.B2(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_211),
.A2(n_222),
.B1(n_228),
.B2(n_227),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_126),
.B(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_214),
.Y(n_272)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_217),
.A2(n_257),
.B1(n_223),
.B2(n_240),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_178),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_218),
.A2(n_256),
.B(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_169),
.A2(n_192),
.B1(n_132),
.B2(n_196),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_132),
.B1(n_192),
.B2(n_122),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_125),
.B(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_125),
.B(n_175),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_237),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_171),
.A2(n_121),
.B(n_125),
.C(n_122),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_179),
.B(n_207),
.C(n_254),
.Y(n_266)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_242),
.Y(n_290)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_125),
.B(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_144),
.B(n_194),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_243),
.B(n_246),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

INVx6_ASAP7_75t_SL g294 ( 
.A(n_244),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_245),
.A2(n_261),
.B1(n_262),
.B2(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_148),
.B(n_194),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_121),
.A2(n_187),
.B(n_162),
.C(n_133),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_218),
.B(n_201),
.C(n_240),
.Y(n_280)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_119),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_255),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_162),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_119),
.B(n_165),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_172),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_149),
.B(n_173),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_266),
.A2(n_300),
.B(n_302),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_270),
.A2(n_244),
.B1(n_282),
.B2(n_301),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_227),
.A2(n_232),
.B1(n_217),
.B2(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_275),
.A2(n_277),
.B1(n_296),
.B2(n_311),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_306),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_207),
.B(n_239),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_292),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_217),
.A2(n_224),
.B1(n_219),
.B2(n_245),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_275),
.B1(n_302),
.B2(n_266),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_208),
.B(n_219),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_287),
.B(n_294),
.C(n_308),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_297),
.C(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_238),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_226),
.A2(n_198),
.B1(n_204),
.B2(n_255),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_SL g297 ( 
.A(n_226),
.B(n_199),
.C(n_247),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_234),
.B(n_251),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_259),
.A2(n_230),
.B1(n_262),
.B2(n_215),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_216),
.A2(n_225),
.B1(n_261),
.B2(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_283),
.B(n_261),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_323),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_279),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_305),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_301),
.B1(n_292),
.B2(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_309),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_326),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_288),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_296),
.A2(n_297),
.B1(n_280),
.B2(n_269),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_324),
.A2(n_333),
.B(n_346),
.Y(n_367)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_280),
.A2(n_287),
.B(n_278),
.C(n_295),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_343),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_273),
.B(n_267),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_268),
.C(n_298),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_339),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_276),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_328),
.B(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_278),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_338),
.Y(n_374)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_295),
.B(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_332),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_311),
.A2(n_291),
.B1(n_265),
.B2(n_263),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_265),
.B(n_307),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_345),
.C(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_264),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_306),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_342),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_294),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_264),
.B(n_293),
.C(n_303),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_281),
.B(n_299),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_274),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_347),
.A2(n_332),
.B(n_342),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_274),
.B(n_291),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_349),
.A2(n_357),
.B(n_359),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_281),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_369),
.C(n_316),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_366),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_320),
.A2(n_310),
.B1(n_303),
.B2(n_299),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_347),
.B1(n_313),
.B2(n_312),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_310),
.B(n_348),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_348),
.B(n_324),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_341),
.A2(n_314),
.B1(n_323),
.B2(n_315),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_362),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_341),
.A2(n_314),
.B1(n_319),
.B2(n_325),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_317),
.A2(n_332),
.B(n_334),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_325),
.B(n_333),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_338),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_339),
.B(n_322),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_356),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_385),
.C(n_369),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_395),
.B1(n_356),
.B2(n_349),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_380),
.A2(n_396),
.B(n_397),
.Y(n_407)
);

AOI22x1_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_336),
.B1(n_331),
.B2(n_329),
.Y(n_381)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_381),
.Y(n_401)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_363),
.B(n_337),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_388),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_318),
.Y(n_384)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_345),
.C(n_328),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_326),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_364),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_390),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_391),
.A2(n_392),
.B1(n_398),
.B2(n_355),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_351),
.A2(n_343),
.B1(n_344),
.B2(n_375),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_373),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_376),
.A2(n_375),
.B1(n_357),
.B2(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_376),
.A2(n_374),
.B1(n_359),
.B2(n_366),
.Y(n_400)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_380),
.A2(n_367),
.B(n_349),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_402),
.A2(n_405),
.B1(n_378),
.B2(n_394),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_406),
.C(n_408),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_350),
.C(n_369),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_360),
.C(n_372),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_388),
.A2(n_374),
.B1(n_353),
.B2(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_410),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_372),
.C(n_367),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_412),
.B(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_396),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_429),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_411),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_427),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_399),
.B1(n_395),
.B2(n_401),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_404),
.B(n_386),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_421),
.B(n_365),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_405),
.A2(n_378),
.B1(n_390),
.B2(n_389),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_420),
.B1(n_401),
.B2(n_418),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_409),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_411),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_415),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_384),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_408),
.C(n_412),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_430),
.B(n_434),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_438),
.B1(n_422),
.B2(n_418),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_416),
.A2(n_407),
.B(n_402),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_414),
.B(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_439),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_407),
.C(n_400),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_429),
.C(n_417),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_443),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_415),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_448),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_425),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_444),
.A2(n_424),
.B1(n_393),
.B2(n_410),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_447),
.Y(n_455)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

OA21x2_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_409),
.B(n_392),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_445),
.A2(n_425),
.B1(n_433),
.B2(n_432),
.Y(n_449)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_446),
.B(n_436),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_454),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_436),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_452),
.A2(n_441),
.B(n_440),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_457),
.A2(n_459),
.B(n_460),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_443),
.C(n_428),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_456),
.A2(n_455),
.B(n_452),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_462),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_449),
.C(n_443),
.Y(n_462)
);

BUFx24_ASAP7_75t_SL g464 ( 
.A(n_463),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_465),
.B(n_458),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_466),
.A2(n_442),
.B(n_393),
.C(n_382),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_453),
.Y(n_468)
);


endmodule