module fake_jpeg_6850_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_22),
.B1(n_15),
.B2(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_18),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_3),
.B(n_4),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_29),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_63),
.Y(n_66)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_17),
.B1(n_36),
.B2(n_26),
.Y(n_70)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_22),
.B1(n_31),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_25),
.B1(n_49),
.B2(n_54),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_62),
.B1(n_51),
.B2(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_29),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_75),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_64),
.B1(n_21),
.B2(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_43),
.B1(n_33),
.B2(n_34),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_80),
.B1(n_52),
.B2(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_82),
.B(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_59),
.B1(n_55),
.B2(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_85),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_94),
.B1(n_101),
.B2(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.C(n_73),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_57),
.C(n_50),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_57),
.B1(n_38),
.B2(n_37),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_119),
.B1(n_38),
.B2(n_18),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_87),
.B1(n_95),
.B2(n_88),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_60),
.A3(n_32),
.B1(n_48),
.B2(n_37),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_48),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_67),
.B1(n_72),
.B2(n_60),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_81),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_88),
.C(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_72),
.C(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_136),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_84),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_129),
.C(n_135),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_94),
.B(n_32),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_131),
.B(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_67),
.B(n_92),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_140),
.B(n_104),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_138),
.B(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_111),
.B1(n_122),
.B2(n_110),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_32),
.C(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_48),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_102),
.B(n_48),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_28),
.B(n_19),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_113),
.B(n_105),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_104),
.C(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_142),
.C(n_129),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_116),
.B(n_28),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_107),
.B1(n_81),
.B2(n_16),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_138),
.B1(n_130),
.B2(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_28),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_153),
.C(n_152),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_124),
.B1(n_128),
.B2(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_16),
.B1(n_13),
.B2(n_5),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_13),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_3),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_142),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_180),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_143),
.C(n_151),
.Y(n_176)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_149),
.C(n_148),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_4),
.Y(n_190)
);

FAx1_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_170),
.CI(n_161),
.CON(n_185),
.SN(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_163),
.B(n_165),
.C(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_158),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_6),
.Y(n_193)
);

OAI21x1_ASAP7_75t_SL g192 ( 
.A1(n_189),
.A2(n_185),
.B(n_186),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_183),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_197),
.B(n_193),
.C(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_194),
.C(n_10),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule