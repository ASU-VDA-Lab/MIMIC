module fake_jpeg_22938_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_16),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_46),
.Y(n_62)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_34),
.Y(n_77)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_58),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_19),
.B1(n_24),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_43),
.B1(n_19),
.B2(n_29),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_71),
.Y(n_94)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_21),
.C(n_34),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_27),
.C(n_26),
.Y(n_109)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_17),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_47),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_32),
.B(n_30),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_88),
.B(n_101),
.C(n_25),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_97),
.B1(n_70),
.B2(n_69),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_98),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_24),
.B(n_47),
.C(n_32),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_47),
.B(n_29),
.C(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_105),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_26),
.B1(n_25),
.B2(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_23),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_72),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_0),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_113),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_127),
.B1(n_105),
.B2(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_130),
.B1(n_85),
.B2(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_71),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_65),
.C(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_57),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_102),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_53),
.B1(n_59),
.B2(n_57),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_102),
.B1(n_104),
.B2(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_53),
.C(n_4),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_109),
.C(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_15),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_86),
.B(n_103),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_142),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_133),
.B1(n_130),
.B2(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_145),
.B1(n_159),
.B2(n_111),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_89),
.C(n_90),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_97),
.B1(n_81),
.B2(n_96),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_90),
.C(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_157),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_99),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_113),
.B(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_99),
.B1(n_98),
.B2(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_162),
.Y(n_177)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_147),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_125),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_180),
.B1(n_154),
.B2(n_161),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_151),
.B(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_117),
.B1(n_116),
.B2(n_119),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_172),
.B1(n_178),
.B2(n_179),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_174),
.C(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_117),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_121),
.B1(n_108),
.B2(n_136),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_134),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_134),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_145),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_127),
.B1(n_7),
.B2(n_9),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_127),
.B1(n_10),
.B2(n_11),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_190),
.C(n_164),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_156),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_183),
.A2(n_188),
.B(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_153),
.A3(n_141),
.B1(n_161),
.B2(n_144),
.C1(n_156),
.C2(n_151),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_196),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_175),
.C(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_190),
.C(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_173),
.B1(n_138),
.B2(n_181),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_210),
.B1(n_189),
.B2(n_173),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_183),
.C(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_218),
.C(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_192),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_186),
.A3(n_185),
.B(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_162),
.C(n_141),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_160),
.C(n_191),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_147),
.B1(n_157),
.B2(n_154),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_202),
.B1(n_209),
.B2(n_155),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_205),
.B(n_198),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_223),
.B(n_227),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_199),
.B(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_211),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_212),
.C(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_199),
.B1(n_159),
.B2(n_150),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_5),
.B(n_10),
.C(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_180),
.Y(n_231)
);

NOR5xp2_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.C(n_223),
.D(n_225),
.E(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_235),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_12),
.B(n_13),
.Y(n_239)
);

AND3x1_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_12),
.C(n_13),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_239),
.B(n_13),
.C(n_14),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_14),
.C(n_15),
.Y(n_241)
);


endmodule