module fake_jpeg_9736_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_19),
.Y(n_63)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_25),
.B(n_29),
.C(n_17),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_22),
.B(n_33),
.C(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_17),
.B1(n_27),
.B2(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_60),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_23),
.B1(n_33),
.B2(n_21),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_19),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_23),
.C(n_33),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_40),
.B(n_34),
.C(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_67),
.B1(n_45),
.B2(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_34),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_13),
.B(n_16),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_90),
.B1(n_75),
.B2(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_77),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_30),
.B(n_18),
.C(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_82),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_20),
.C(n_8),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_48),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

OR2x6_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_44),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_62),
.A3(n_34),
.B1(n_20),
.B2(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_65),
.B1(n_68),
.B2(n_83),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_90),
.B1(n_91),
.B2(n_65),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_119),
.B1(n_66),
.B2(n_78),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.C(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_64),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_64),
.C(n_20),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_34),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_8),
.B1(n_14),
.B2(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_124),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_125),
.B(n_132),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_134),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_128),
.B(n_137),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_85),
.B(n_92),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_99),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_94),
.B1(n_102),
.B2(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_82),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_79),
.B(n_72),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_103),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_69),
.B1(n_81),
.B2(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_74),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_100),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_77),
.B1(n_88),
.B2(n_74),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_88),
.B1(n_86),
.B2(n_3),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_9),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_113),
.C(n_94),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_86),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_9),
.B1(n_14),
.B2(n_4),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_149),
.B1(n_102),
.B2(n_107),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_150),
.A2(n_157),
.B(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_155),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_159),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_106),
.A3(n_101),
.B1(n_99),
.B2(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_106),
.B1(n_97),
.B2(n_101),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_122),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_161),
.C(n_174),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_170),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_167),
.B(n_2),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_173),
.B(n_4),
.Y(n_201)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_1),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_143),
.B(n_127),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_198),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_145),
.B1(n_133),
.B2(n_141),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_193),
.B1(n_190),
.B2(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_130),
.C(n_146),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_140),
.C(n_134),
.Y(n_188)
);

AOI21x1_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_128),
.B(n_149),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_137),
.C(n_121),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_192),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_148),
.B1(n_2),
.B2(n_1),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_9),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_163),
.B1(n_167),
.B2(n_153),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_215),
.B(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_166),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_161),
.C(n_154),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_173),
.B1(n_156),
.B2(n_178),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_201),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_156),
.B1(n_162),
.B2(n_151),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_183),
.B1(n_189),
.B2(n_193),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_150),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_189),
.B(n_195),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_171),
.B1(n_150),
.B2(n_7),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_179),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_227),
.C(n_232),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_179),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_196),
.B1(n_192),
.B2(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

AOI31xp67_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_187),
.A3(n_200),
.B(n_191),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_233),
.B(n_237),
.C(n_239),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_185),
.C(n_188),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_207),
.B1(n_215),
.B2(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_206),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_194),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_240),
.B(n_242),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_245),
.B1(n_234),
.B2(n_235),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_209),
.B1(n_203),
.B2(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_220),
.B1(n_219),
.B2(n_210),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_214),
.B(n_204),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_5),
.C(n_6),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_249),
.B(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_7),
.C(n_11),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_226),
.B1(n_230),
.B2(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_237),
.B1(n_226),
.B2(n_224),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_244),
.B(n_242),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_259),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_255),
.B(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_267),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_R g267 ( 
.A(n_255),
.B(n_248),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_253),
.B(n_244),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_272),
.B(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_11),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_275),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_276),
.A2(n_12),
.B1(n_15),
.B2(n_274),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_12),
.B(n_15),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_277),
.Y(n_280)
);


endmodule