module real_aes_7112_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_0), .A2(n_7), .B1(n_441), .B2(n_712), .C1(n_717), .C2(n_718), .Y(n_440) );
INVx1_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_2), .A2(n_142), .B(n_147), .C(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_3), .A2(n_137), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g453 ( .A(n_4), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_5), .B(n_161), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_6), .B(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_7), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_8), .A2(n_137), .B(n_471), .Y(n_470) );
AND2x6_ASAP7_75t_L g142 ( .A(n_9), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g171 ( .A(n_10), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_11), .B(n_43), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_11), .B(n_43), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_12), .A2(n_249), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_13), .B(n_152), .Y(n_188) );
INVx1_ASAP7_75t_L g475 ( .A(n_14), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_15), .B(n_151), .Y(n_523) );
INVx1_ASAP7_75t_L g135 ( .A(n_16), .Y(n_135) );
INVx1_ASAP7_75t_L g535 ( .A(n_17), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_18), .A2(n_172), .B(n_197), .C(n_199), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_19), .B(n_161), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_20), .B(n_464), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_21), .B(n_137), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_22), .B(n_257), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_23), .A2(n_151), .B(n_153), .C(n_157), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_24), .B(n_161), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_25), .B(n_152), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_26), .A2(n_155), .B(n_199), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_27), .B(n_152), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_28), .Y(n_217) );
INVx1_ASAP7_75t_L g231 ( .A(n_29), .Y(n_231) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_30), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_31), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_32), .B(n_152), .Y(n_454) );
INVx1_ASAP7_75t_L g254 ( .A(n_33), .Y(n_254) );
INVx1_ASAP7_75t_L g488 ( .A(n_34), .Y(n_488) );
INVx2_ASAP7_75t_L g140 ( .A(n_35), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_36), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_37), .A2(n_151), .B(n_210), .C(n_212), .Y(n_209) );
INVxp67_ASAP7_75t_L g255 ( .A(n_38), .Y(n_255) );
CKINVDCx14_ASAP7_75t_R g208 ( .A(n_39), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_40), .A2(n_147), .B(n_230), .C(n_236), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_41), .A2(n_142), .B(n_147), .C(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_42), .A2(n_120), .B1(n_121), .B2(n_428), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_42), .Y(n_428) );
INVx1_ASAP7_75t_L g487 ( .A(n_44), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_45), .A2(n_169), .B(n_170), .C(n_173), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_46), .B(n_152), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_47), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_48), .Y(n_251) );
INVx1_ASAP7_75t_L g145 ( .A(n_49), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_50), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_51), .B(n_137), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_52), .A2(n_147), .B1(n_157), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_53), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_54), .Y(n_450) );
CKINVDCx14_ASAP7_75t_R g167 ( .A(n_55), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_56), .A2(n_169), .B(n_212), .C(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_57), .Y(n_516) );
INVx1_ASAP7_75t_L g472 ( .A(n_58), .Y(n_472) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
INVx1_ASAP7_75t_L g134 ( .A(n_60), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_61), .A2(n_100), .B1(n_113), .B2(n_723), .Y(n_99) );
INVx1_ASAP7_75t_SL g211 ( .A(n_62), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_63), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_64), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g220 ( .A(n_65), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_66), .A2(n_212), .B(n_464), .C(n_465), .Y(n_463) );
INVxp67_ASAP7_75t_L g466 ( .A(n_67), .Y(n_466) );
INVx1_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_69), .A2(n_137), .B(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_70), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_71), .A2(n_137), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_72), .Y(n_491) );
INVx1_ASAP7_75t_L g510 ( .A(n_73), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_74), .A2(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g195 ( .A(n_75), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_76), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_77), .A2(n_142), .B(n_147), .C(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_78), .A2(n_137), .B(n_144), .Y(n_136) );
INVx1_ASAP7_75t_L g198 ( .A(n_79), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_80), .B(n_232), .Y(n_504) );
INVx2_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g185 ( .A(n_82), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_83), .B(n_464), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_84), .A2(n_142), .B(n_147), .C(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g109 ( .A(n_85), .Y(n_109) );
OR2x2_ASAP7_75t_L g432 ( .A(n_85), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g711 ( .A(n_85), .B(n_434), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_86), .A2(n_147), .B(n_219), .C(n_222), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_87), .B(n_164), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_88), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_89), .A2(n_142), .B(n_147), .C(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_90), .Y(n_527) );
INVx1_ASAP7_75t_L g462 ( .A(n_91), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_92), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_93), .B(n_232), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_94), .B(n_130), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_95), .B(n_130), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_98), .A2(n_137), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g723 ( .A(n_102), .Y(n_723) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g434 ( .A(n_108), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g710 ( .A(n_109), .B(n_434), .Y(n_710) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_109), .B(n_433), .Y(n_720) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_439), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g722 ( .A(n_117), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_429), .B(n_436), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_122), .A2(n_442), .B1(n_710), .B2(n_711), .Y(n_441) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g716 ( .A(n_123), .Y(n_716) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_354), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_296), .C(n_326), .D(n_336), .Y(n_124) );
OAI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_201), .B(n_259), .C(n_286), .Y(n_125) );
OAI222xp33_ASAP7_75t_L g381 ( .A1(n_126), .A2(n_301), .B1(n_382), .B2(n_383), .C1(n_384), .C2(n_385), .Y(n_381) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_176), .Y(n_126) );
AOI33xp33_ASAP7_75t_L g307 ( .A1(n_127), .A2(n_294), .A3(n_295), .B1(n_308), .B2(n_313), .B3(n_315), .Y(n_307) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_127), .A2(n_365), .B(n_367), .C(n_369), .Y(n_364) );
OR2x2_ASAP7_75t_L g380 ( .A(n_127), .B(n_366), .Y(n_380) );
INVx1_ASAP7_75t_L g413 ( .A(n_127), .Y(n_413) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
INVx2_ASAP7_75t_L g290 ( .A(n_128), .Y(n_290) );
AND2x2_ASAP7_75t_L g306 ( .A(n_128), .B(n_192), .Y(n_306) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_128), .Y(n_341) );
AND2x2_ASAP7_75t_L g370 ( .A(n_128), .B(n_163), .Y(n_370) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_160), .Y(n_128) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_129), .A2(n_193), .B(n_200), .Y(n_192) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_129), .A2(n_206), .B(n_214), .Y(n_205) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_130), .A2(n_460), .B(n_467), .Y(n_459) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g247 ( .A(n_131), .Y(n_247) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_132), .B(n_133), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx2_ASAP7_75t_L g249 ( .A(n_137), .Y(n_249) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_138), .B(n_142), .Y(n_182) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g235 ( .A(n_139), .Y(n_235) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
INVx1_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
INVx3_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
INVx1_ASAP7_75t_L g464 ( .A(n_141), .Y(n_464) );
INVx4_ASAP7_75t_SL g159 ( .A(n_142), .Y(n_159) );
BUFx3_ASAP7_75t_L g236 ( .A(n_142), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_159), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_SL g166 ( .A1(n_146), .A2(n_159), .B(n_167), .C(n_168), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_146), .A2(n_159), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_146), .A2(n_159), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_146), .A2(n_159), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_146), .A2(n_159), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_146), .A2(n_159), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_146), .A2(n_159), .B(n_532), .C(n_533), .Y(n_531) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_151), .B(n_211), .Y(n_210) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_155), .B(n_198), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_155), .A2(n_232), .B1(n_254), .B2(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_155), .B(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_156), .A2(n_187), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g455 ( .A(n_157), .Y(n_455) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_159), .A2(n_182), .B1(n_485), .B2(n_489), .Y(n_484) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_161), .A2(n_470), .B(n_476), .Y(n_469) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_162), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_162), .A2(n_216), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_162), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g506 ( .A(n_162), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g270 ( .A(n_163), .Y(n_270) );
BUFx3_ASAP7_75t_L g278 ( .A(n_163), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_163), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g289 ( .A(n_163), .B(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_163), .B(n_177), .Y(n_318) );
AND2x2_ASAP7_75t_L g387 ( .A(n_163), .B(n_321), .Y(n_387) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_175), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx2_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_164), .A2(n_182), .B(n_228), .C(n_229), .Y(n_227) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_164), .A2(n_530), .B(n_536), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx5_ASAP7_75t_L g232 ( .A(n_172), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_172), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_172), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g189 ( .A(n_173), .Y(n_189) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g199 ( .A(n_174), .Y(n_199) );
INVx2_ASAP7_75t_SL g281 ( .A(n_176), .Y(n_281) );
OR2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_177), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g323 ( .A(n_177), .Y(n_323) );
AND2x2_ASAP7_75t_L g334 ( .A(n_177), .B(n_290), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_177), .B(n_319), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_177), .B(n_321), .Y(n_366) );
AND2x2_ASAP7_75t_L g425 ( .A(n_177), .B(n_370), .Y(n_425) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g295 ( .A(n_178), .B(n_192), .Y(n_295) );
AND2x2_ASAP7_75t_L g305 ( .A(n_178), .B(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g327 ( .A(n_178), .Y(n_327) );
AND3x2_ASAP7_75t_L g386 ( .A(n_178), .B(n_387), .C(n_388), .Y(n_386) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_190), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_179), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_179), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_179), .B(n_527), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_182), .A2(n_217), .B(n_218), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_182), .A2(n_450), .B(n_451), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_182), .A2(n_510), .B(n_511), .Y(n_509) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_189), .B(n_220), .C(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_189), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_189), .A2(n_513), .B(n_514), .Y(n_512) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_192), .Y(n_277) );
INVx1_ASAP7_75t_SL g321 ( .A(n_192), .Y(n_321) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_192), .B(n_270), .C(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_239), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_202), .A2(n_305), .B(n_357), .C(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_204), .B(n_226), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_204), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g373 ( .A(n_204), .Y(n_373) );
AND2x2_ASAP7_75t_L g394 ( .A(n_204), .B(n_241), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_204), .B(n_303), .Y(n_422) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
AND2x2_ASAP7_75t_L g267 ( .A(n_205), .B(n_258), .Y(n_267) );
INVx2_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
AND2x2_ASAP7_75t_L g294 ( .A(n_205), .B(n_241), .Y(n_294) );
AND2x2_ASAP7_75t_L g344 ( .A(n_205), .B(n_226), .Y(n_344) );
INVx1_ASAP7_75t_L g348 ( .A(n_205), .Y(n_348) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_213), .Y(n_524) );
INVx2_ASAP7_75t_SL g258 ( .A(n_215), .Y(n_258) );
BUFx2_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
AND2x2_ASAP7_75t_L g411 ( .A(n_215), .B(n_226), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx1_ASAP7_75t_L g257 ( .A(n_225), .Y(n_257) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_225), .A2(n_519), .B(n_526), .Y(n_518) );
INVx3_ASAP7_75t_SL g241 ( .A(n_226), .Y(n_241) );
AND2x2_ASAP7_75t_L g266 ( .A(n_226), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g273 ( .A(n_226), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g303 ( .A(n_226), .B(n_263), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_226), .B(n_258), .Y(n_312) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_226), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_226), .B(n_288), .Y(n_335) );
AND2x2_ASAP7_75t_L g363 ( .A(n_226), .B(n_243), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_226), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_226), .B(n_242), .Y(n_401) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_237), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .C(n_234), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_232), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_235), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x2_ASAP7_75t_L g325 ( .A(n_241), .B(n_274), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_241), .B(n_267), .Y(n_353) );
AND2x2_ASAP7_75t_L g371 ( .A(n_241), .B(n_288), .Y(n_371) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_258), .Y(n_242) );
AND2x2_ASAP7_75t_L g272 ( .A(n_243), .B(n_258), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_243), .B(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g310 ( .A(n_243), .Y(n_310) );
OR2x2_ASAP7_75t_L g358 ( .A(n_243), .B(n_278), .Y(n_358) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .B(n_256), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_245), .A2(n_264), .B(n_265), .Y(n_263) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_245), .A2(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_SL g500 ( .A1(n_246), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_247), .A2(n_449), .B(n_456), .Y(n_448) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_247), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_247), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g264 ( .A(n_248), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_256), .Y(n_265) );
AND2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_263), .Y(n_293) );
INVx1_ASAP7_75t_L g301 ( .A(n_258), .Y(n_301) );
AND2x2_ASAP7_75t_L g396 ( .A(n_258), .B(n_274), .Y(n_396) );
AOI222xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_268), .B1(n_271), .B2(n_275), .C1(n_279), .C2(n_282), .Y(n_259) );
INVx1_ASAP7_75t_L g391 ( .A(n_260), .Y(n_391) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_266), .Y(n_260) );
AND2x2_ASAP7_75t_L g287 ( .A(n_261), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g298 ( .A(n_261), .B(n_267), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_261), .B(n_289), .Y(n_314) );
OAI222xp33_ASAP7_75t_L g336 ( .A1(n_261), .A2(n_337), .B1(n_342), .B2(n_343), .C1(n_351), .C2(n_353), .Y(n_336) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g324 ( .A(n_263), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_263), .B(n_344), .Y(n_384) );
AND2x2_ASAP7_75t_L g395 ( .A(n_263), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g403 ( .A(n_266), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_268), .B(n_319), .Y(n_382) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_270), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g340 ( .A(n_270), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx3_ASAP7_75t_L g285 ( .A(n_273), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g375 ( .A1(n_273), .A2(n_376), .B(n_379), .C(n_381), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_273), .B(n_310), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_273), .B(n_293), .Y(n_415) );
AND2x2_ASAP7_75t_L g288 ( .A(n_274), .B(n_284), .Y(n_288) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_278), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g367 ( .A(n_278), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g406 ( .A(n_278), .B(n_306), .Y(n_406) );
INVx1_ASAP7_75t_L g418 ( .A(n_278), .Y(n_418) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_281), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g399 ( .A(n_284), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B(n_291), .C(n_295), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_287), .A2(n_317), .B1(n_332), .B2(n_335), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_288), .B(n_302), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_288), .B(n_310), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_289), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g352 ( .A(n_289), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_289), .B(n_339), .Y(n_359) );
INVx2_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NOR4xp25_ASAP7_75t_L g297 ( .A(n_294), .B(n_298), .C(n_299), .D(n_302), .Y(n_297) );
INVx1_ASAP7_75t_SL g368 ( .A(n_295), .Y(n_368) );
AND2x2_ASAP7_75t_L g412 ( .A(n_295), .B(n_413), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_304), .B(n_307), .C(n_316), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_303), .B(n_373), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_305), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_SL g378 ( .A(n_306), .Y(n_378) );
AND2x2_ASAP7_75t_L g417 ( .A(n_306), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_310), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_314), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_315), .B(n_340), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_322), .B(n_324), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g392 ( .A(n_319), .Y(n_392) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_L g420 ( .A(n_320), .Y(n_420) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B(n_331), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_327), .Y(n_339) );
OR2x2_ASAP7_75t_L g377 ( .A(n_327), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_330), .A2(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_334), .A2(n_361), .B1(n_364), .B2(n_371), .C(n_372), .Y(n_360) );
INVx1_ASAP7_75t_SL g404 ( .A(n_335), .Y(n_404) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g351 ( .A(n_339), .B(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B1(n_348), .B2(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_347), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR4xp25_ASAP7_75t_L g354 ( .A(n_355), .B(n_389), .C(n_402), .D(n_414), .Y(n_354) );
NAND3xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_360), .C(n_375), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_358), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_365), .B(n_370), .Y(n_374) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_377), .A2(n_403), .B1(n_404), .B2(n_405), .C(n_407), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_379), .A2(n_394), .B(n_395), .C(n_397), .Y(n_393) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_380), .A2(n_398), .B1(n_400), .B2(n_401), .Y(n_397) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_392), .C(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g408 ( .A(n_401), .Y(n_408) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_409), .B(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B1(n_419), .B2(n_421), .C(n_423), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_432), .Y(n_438) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_436), .A2(n_440), .B(n_721), .Y(n_439) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g713 ( .A(n_442), .Y(n_713) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_626), .Y(n_442) );
NOR5xp2_ASAP7_75t_L g443 ( .A(n_444), .B(n_549), .C(n_581), .D(n_596), .E(n_613), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_477), .B(n_496), .C(n_537), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_458), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_446), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_446), .B(n_601), .Y(n_664) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_447), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_447), .B(n_493), .Y(n_550) );
AND2x2_ASAP7_75t_L g591 ( .A(n_447), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_447), .B(n_560), .Y(n_595) );
OR2x2_ASAP7_75t_L g632 ( .A(n_447), .B(n_483), .Y(n_632) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g482 ( .A(n_448), .B(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g540 ( .A(n_448), .Y(n_540) );
OR2x2_ASAP7_75t_L g703 ( .A(n_448), .B(n_543), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_458), .A2(n_606), .B1(n_607), .B2(n_610), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_458), .B(n_540), .Y(n_689) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .Y(n_458) );
AND2x2_ASAP7_75t_L g495 ( .A(n_459), .B(n_483), .Y(n_495) );
AND2x2_ASAP7_75t_L g542 ( .A(n_459), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g547 ( .A(n_459), .Y(n_547) );
INVx3_ASAP7_75t_L g560 ( .A(n_459), .Y(n_560) );
OR2x2_ASAP7_75t_L g580 ( .A(n_459), .B(n_543), .Y(n_580) );
AND2x2_ASAP7_75t_L g599 ( .A(n_459), .B(n_469), .Y(n_599) );
BUFx2_ASAP7_75t_L g631 ( .A(n_459), .Y(n_631) );
AND2x4_ASAP7_75t_L g546 ( .A(n_468), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g481 ( .A(n_469), .Y(n_481) );
INVx2_ASAP7_75t_L g494 ( .A(n_469), .Y(n_494) );
OR2x2_ASAP7_75t_L g562 ( .A(n_469), .B(n_543), .Y(n_562) );
AND2x2_ASAP7_75t_L g592 ( .A(n_469), .B(n_483), .Y(n_592) );
AND2x2_ASAP7_75t_L g609 ( .A(n_469), .B(n_540), .Y(n_609) );
AND2x2_ASAP7_75t_L g649 ( .A(n_469), .B(n_560), .Y(n_649) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_469), .B(n_495), .Y(n_685) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp33_ASAP7_75t_SL g478 ( .A(n_479), .B(n_492), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_480), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_481), .A2(n_495), .B(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_481), .B(n_483), .Y(n_679) );
AND2x2_ASAP7_75t_L g615 ( .A(n_482), .B(n_616), .Y(n_615) );
INVx3_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_483), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_492), .B(n_540), .Y(n_708) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_493), .A2(n_651), .B1(n_652), .B2(n_657), .Y(n_650) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g579 ( .A(n_494), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g616 ( .A(n_494), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_495), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g670 ( .A(n_495), .Y(n_670) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_517), .Y(n_497) );
INVx4_ASAP7_75t_L g556 ( .A(n_498), .Y(n_556) );
AND2x2_ASAP7_75t_L g634 ( .A(n_498), .B(n_601), .Y(n_634) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx3_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
AND2x2_ASAP7_75t_L g567 ( .A(n_499), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
INVx2_ASAP7_75t_L g585 ( .A(n_499), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_499), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g642 ( .A(n_499), .B(n_637), .Y(n_642) );
AND2x2_ASAP7_75t_L g707 ( .A(n_499), .B(n_677), .Y(n_707) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g548 ( .A(n_508), .B(n_529), .Y(n_548) );
INVx2_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g619 ( .A(n_517), .B(n_567), .Y(n_619) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx2_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
INVx1_ASAP7_75t_L g566 ( .A(n_518), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_518), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_518), .B(n_568), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
AND2x2_ASAP7_75t_L g601 ( .A(n_528), .B(n_558), .Y(n_601) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g554 ( .A(n_529), .Y(n_554) );
AND2x2_ASAP7_75t_L g637 ( .A(n_529), .B(n_568), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_544), .B(n_548), .Y(n_537) );
INVx1_ASAP7_75t_SL g582 ( .A(n_538), .Y(n_582) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_539), .B(n_546), .Y(n_639) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g588 ( .A(n_540), .B(n_543), .Y(n_588) );
AND2x2_ASAP7_75t_L g617 ( .A(n_540), .B(n_561), .Y(n_617) );
OR2x2_ASAP7_75t_L g620 ( .A(n_540), .B(n_580), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_541), .A2(n_633), .B1(n_685), .B2(n_686), .C1(n_688), .C2(n_690), .Y(n_684) );
BUFx2_ASAP7_75t_L g598 ( .A(n_543), .Y(n_598) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g587 ( .A(n_546), .B(n_588), .Y(n_587) );
INVx3_ASAP7_75t_SL g604 ( .A(n_546), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_546), .B(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g593 ( .A(n_548), .B(n_553), .Y(n_593) );
INVx1_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_551), .B1(n_555), .B2(n_559), .C(n_563), .Y(n_549) );
OR2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g606 ( .A(n_553), .B(n_576), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_553), .B(n_566), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_553), .B(n_601), .Y(n_651) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_553), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g672 ( .A(n_553), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g557 ( .A(n_554), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_554), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_554), .B(n_572), .Y(n_603) );
INVx1_ASAP7_75t_L g669 ( .A(n_554), .Y(n_669) );
INVx1_ASAP7_75t_L g644 ( .A(n_555), .Y(n_644) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g656 ( .A(n_556), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g668 ( .A(n_556), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g673 ( .A(n_557), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_557), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g576 ( .A(n_558), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_558), .B(n_568), .Y(n_589) );
INVx1_ASAP7_75t_L g655 ( .A(n_558), .Y(n_655) );
INVx1_ASAP7_75t_L g676 ( .A(n_559), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI21xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_569), .B(n_578), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g709 ( .A(n_565), .B(n_642), .Y(n_709) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g677 ( .A(n_566), .B(n_637), .Y(n_677) );
AOI32xp33_ASAP7_75t_L g590 ( .A1(n_567), .A2(n_573), .A3(n_591), .B1(n_593), .B2(n_594), .Y(n_590) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_567), .A2(n_599), .A3(n_682), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_697), .Y(n_692) );
INVx2_ASAP7_75t_L g572 ( .A(n_568), .Y(n_572) );
INVx1_ASAP7_75t_L g682 ( .A(n_568), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_570), .B(n_576), .Y(n_625) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_571), .B(n_637), .Y(n_687) );
INVx1_ASAP7_75t_L g574 ( .A(n_572), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_572), .B(n_601), .Y(n_691) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_580), .B(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_583), .B1(n_586), .B2(n_589), .C(n_590), .Y(n_581) );
OR2x2_ASAP7_75t_L g602 ( .A(n_583), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g611 ( .A(n_583), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g636 ( .A(n_584), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g640 ( .A(n_594), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B1(n_602), .B2(n_604), .C(n_605), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_598), .A2(n_629), .B1(n_633), .B2(n_634), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_599), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_599), .Y(n_704) );
INVx1_ASAP7_75t_L g698 ( .A(n_601), .Y(n_698) );
INVx1_ASAP7_75t_SL g633 ( .A(n_602), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_604), .B(n_632), .Y(n_694) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_609), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g675 ( .A(n_609), .Y(n_675) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_618), .B1(n_620), .B2(n_621), .C(n_623), .Y(n_613) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_615), .A2(n_633), .B1(n_679), .B2(n_680), .Y(n_678) );
CKINVDCx14_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_620), .A2(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_659), .C(n_683), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_635), .C(n_643), .D(n_650), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g706 ( .A(n_631), .Y(n_706) );
INVx3_ASAP7_75t_SL g700 ( .A(n_632), .Y(n_700) );
OR2x2_ASAP7_75t_L g705 ( .A(n_632), .B(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B1(n_640), .B2(n_642), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_637), .B(n_655), .Y(n_696) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B(n_647), .Y(n_643) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_662), .B(n_665), .C(n_678), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g693 ( .A(n_664), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B1(n_671), .B2(n_674), .C1(n_676), .C2(n_677), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_675), .B(n_703), .C(n_704), .D(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_692), .C(n_701), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_710), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_711), .Y(n_715) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
endmodule