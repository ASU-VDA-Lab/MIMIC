module real_jpeg_2517_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_64),
.B1(n_67),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_24),
.C(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_2),
.B(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_37),
.B1(n_64),
.B2(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_2),
.B(n_44),
.C(n_48),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_62),
.C(n_64),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_55),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_78),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_137),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_30),
.B1(n_64),
.B2(n_67),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_9),
.A2(n_52),
.B1(n_64),
.B2(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_52),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_16),
.B(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.C(n_86),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_17),
.A2(n_18),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_19),
.B(n_40),
.C(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_27),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_25),
.B(n_132),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_28),
.B(n_34),
.Y(n_110)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_53),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_42),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_70)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_48),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_54),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21x1_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_68),
.B(n_71),
.Y(n_58)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_60),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_64),
.B(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_69),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_69),
.B(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_72),
.B(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_86),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_84),
.B2(n_85),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_84),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B(n_81),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_82),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_77),
.A2(n_83),
.B(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_77),
.B(n_172),
.Y(n_186)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_78),
.B(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_83),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_81),
.B(n_185),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_92),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_95),
.B(n_186),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_98),
.B(n_171),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_113),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_112),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_105),
.B(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_138),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_143),
.B(n_204),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_140),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_134),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_126),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_134),
.B1(n_135),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21x1_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_158),
.B(n_203),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_156),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_198),
.B(n_202),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_180),
.B(n_197),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_173),
.B1(n_174),
.B2(n_179),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_187),
.B(n_196),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_184),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B(n_195),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);


endmodule