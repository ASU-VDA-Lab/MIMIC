module real_jpeg_13362_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.C(n_27),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_2),
.B(n_74),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_35),
.C(n_49),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g106 ( 
.A(n_2),
.B(n_60),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_2),
.A2(n_80),
.B(n_112),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_46),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_90)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_94),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_64),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_17),
.B(n_64),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.C(n_55),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_18),
.B(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_30),
.Y(n_85)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_20),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_20),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_23),
.B(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_23),
.B(n_31),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_24),
.A2(n_25),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_28),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B(n_39),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_31),
.A2(n_33),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_31),
.A2(n_39),
.B(n_117),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_32),
.B(n_41),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_32),
.A2(n_40),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_34),
.B(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_43),
.A2(n_55),
.B1(n_56),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_43),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_51),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_47),
.B(n_90),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_63),
.Y(n_70)
);

NOR2x1_ASAP7_75t_R g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_83),
.B2(n_84),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_89),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_132),
.B(n_137),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_113),
.B(n_131),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_121),
.B(n_130),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_119),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_125),
.B(n_129),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);


endmodule