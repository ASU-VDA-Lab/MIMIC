module fake_jpeg_10705_n_219 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_31),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_8),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_48),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_20),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_24),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_42),
.B1(n_41),
.B2(n_25),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_98),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_31),
.B(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_27),
.B1(n_24),
.B2(n_28),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_105),
.B1(n_73),
.B2(n_65),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_104),
.B1(n_66),
.B2(n_62),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_36),
.C(n_29),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_60),
.C(n_35),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_26),
.B1(n_35),
.B2(n_47),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_55),
.B(n_74),
.C(n_77),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_35),
.B(n_3),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_95),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_11),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_128),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_12),
.C(n_15),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.C(n_4),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_62),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_15),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_90),
.B1(n_82),
.B2(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_136),
.B1(n_149),
.B2(n_119),
.Y(n_153)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_85),
.B1(n_81),
.B2(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_142),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_83),
.B1(n_95),
.B2(n_106),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_107),
.B1(n_118),
.B2(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_2),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_3),
.B(n_4),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_121),
.B(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_6),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_162),
.B1(n_169),
.B2(n_140),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_123),
.B1(n_115),
.B2(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_111),
.B(n_121),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_146),
.B(n_144),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

NOR2x1_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_149),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_133),
.C(n_145),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_180),
.C(n_162),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_132),
.Y(n_180)
);

AO21x2_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_130),
.B(n_133),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_181),
.A2(n_182),
.B1(n_169),
.B2(n_168),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_180),
.C(n_182),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_151),
.B(n_131),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_190),
.B(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_143),
.Y(n_187)
);

AOI31xp67_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_191),
.A3(n_177),
.B(n_176),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_171),
.B1(n_181),
.B2(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_151),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_153),
.B1(n_165),
.B2(n_152),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_176),
.Y(n_201)
);

AOI21x1_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_172),
.B(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_192),
.B(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_198),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_181),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_202),
.B1(n_181),
.B2(n_193),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_198),
.B(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_188),
.B1(n_160),
.B2(n_163),
.Y(n_206)
);

NAND4xp25_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.C(n_161),
.D(n_107),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_203),
.B(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_208),
.C(n_209),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_216),
.B(n_213),
.Y(n_219)
);


endmodule