module fake_netlist_1_11496_n_286 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_286);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_286;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_214;
wire n_267;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_244;
wire n_102;
wire n_141;
wire n_119;
wire n_115;
wire n_97;
wire n_167;
wire n_284;
wire n_107;
wire n_158;
wire n_278;
wire n_114;
wire n_121;
wire n_94;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_254;
wire n_161;
wire n_262;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_180;
wire n_104;
wire n_277;
wire n_160;
wire n_98;
wire n_276;
wire n_154;
wire n_272;
wire n_285;
wire n_195;
wire n_165;
wire n_146;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_215;
wire n_155;
wire n_116;
wire n_108;
wire n_209;
wire n_217;
wire n_139;
wire n_229;
wire n_230;
wire n_274;
wire n_198;
wire n_169;
wire n_193;
wire n_273;
wire n_282;
wire n_252;
wire n_152;
wire n_113;
wire n_241;
wire n_156;
wire n_95;
wire n_124;
wire n_238;
wire n_128;
wire n_129;
wire n_120;
wire n_206;
wire n_245;
wire n_135;
wire n_188;
wire n_201;
wire n_197;
wire n_242;
wire n_260;
wire n_247;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_202;
wire n_210;
wire n_142;
wire n_184;
wire n_265;
wire n_191;
wire n_264;
wire n_281;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_275;
wire n_178;
wire n_118;
wire n_258;
wire n_253;
wire n_179;
wire n_131;
wire n_112;
wire n_266;
wire n_205;
wire n_143;
wire n_213;
wire n_243;
wire n_235;
wire n_182;
wire n_263;
wire n_166;
wire n_162;
wire n_186;
wire n_163;
wire n_226;
wire n_174;
wire n_159;
wire n_105;
wire n_227;
wire n_268;
wire n_248;
wire n_231;
wire n_136;
wire n_283;
wire n_176;
wire n_144;
wire n_183;
wire n_256;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_261;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_271;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_270;
wire n_246;
wire n_153;
wire n_259;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_93;
wire n_151;
wire n_140;
wire n_207;
wire n_257;
wire n_224;
wire n_96;
wire n_269;
wire n_225;
wire n_279;
BUFx2_ASAP7_75t_L g92 ( .A(n_79), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_37), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_47), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_45), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_16), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_68), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_85), .B(n_91), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_66), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_80), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_60), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_40), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_82), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_12), .Y(n_113) );
BUFx5_ASAP7_75t_L g114 ( .A(n_35), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_24), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_26), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_29), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_53), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_89), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_14), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_46), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_56), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_55), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_42), .Y(n_130) );
BUFx10_ASAP7_75t_L g131 ( .A(n_22), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_62), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_73), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_77), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_44), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_63), .Y(n_136) );
BUFx10_ASAP7_75t_L g137 ( .A(n_34), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_23), .Y(n_138) );
INVx2_ASAP7_75t_SL g139 ( .A(n_18), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_11), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_114), .B(n_13), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_92), .B(n_0), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_127), .B(n_0), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_131), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_111), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_134), .B(n_1), .Y(n_151) );
AOI22xp33_ASAP7_75t_SL g152 ( .A1(n_140), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_137), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_137), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_94), .B(n_2), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_139), .B(n_4), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_99), .Y(n_162) );
AOI22xp33_ASAP7_75t_SL g163 ( .A1(n_113), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_163) );
BUFx10_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_141), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVxp67_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_155), .B(n_109), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_147), .B(n_129), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_159), .B(n_114), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_156), .B(n_130), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_161), .B(n_114), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_168), .B(n_146), .Y(n_179) );
BUFx5_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_173), .B(n_143), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_173), .B(n_144), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_164), .B(n_161), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_176), .A2(n_145), .B(n_149), .C(n_128), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_164), .B(n_149), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_165), .B(n_95), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_166), .B(n_152), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_178), .A2(n_132), .B1(n_112), .B2(n_163), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_171), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_172), .B(n_103), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_177), .B(n_106), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_179), .B(n_177), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_190), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_187), .A2(n_178), .B1(n_174), .B2(n_142), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_183), .A2(n_174), .B(n_101), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_181), .B(n_116), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_180), .A2(n_96), .B1(n_97), .B2(n_93), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_184), .A2(n_100), .B(n_102), .C(n_98), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_180), .B(n_104), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_186), .A2(n_108), .B(n_105), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_189), .A2(n_117), .B1(n_110), .B2(n_115), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_188), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_201), .A2(n_196), .B(n_193), .Y(n_205) );
AO22x2_ASAP7_75t_L g206 ( .A1(n_203), .A2(n_192), .B1(n_191), .B2(n_185), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_204), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_200), .A2(n_123), .B(n_120), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_195), .A2(n_138), .B1(n_119), .B2(n_122), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_198), .B(n_124), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_202), .A2(n_126), .B(n_125), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_197), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_194), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_199), .B(n_133), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_212), .B(n_8), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_207), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_210), .B(n_9), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_210), .B(n_135), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_213), .Y(n_219) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_205), .A2(n_121), .B(n_148), .Y(n_220) );
AOI21x1_ASAP7_75t_L g221 ( .A1(n_206), .A2(n_154), .B(n_150), .Y(n_221) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_208), .A2(n_157), .B(n_160), .Y(n_222) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_214), .A2(n_158), .A3(n_175), .B(n_170), .Y(n_223) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_211), .A2(n_158), .B(n_175), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_207), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_15), .B(n_17), .Y(n_228) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_19), .A3(n_20), .B(n_21), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_226), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_220), .A2(n_27), .B(n_28), .Y(n_231) );
OR2x6_ASAP7_75t_L g232 ( .A(n_215), .B(n_30), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_217), .B(n_31), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_216), .Y(n_234) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_221), .A2(n_32), .B(n_33), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_227), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_224), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_224), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_36), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_225), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
INVxp67_ASAP7_75t_SL g242 ( .A(n_222), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_229), .B(n_39), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_219), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_230), .B(n_48), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_245), .B(n_49), .Y(n_247) );
AOI21x1_ASAP7_75t_L g248 ( .A1(n_238), .A2(n_54), .B(n_57), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_232), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_234), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_236), .B(n_90), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_233), .B(n_59), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_240), .B(n_61), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_64), .B(n_65), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_239), .B(n_67), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_244), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_256) );
AOI211xp5_ASAP7_75t_SL g257 ( .A1(n_243), .A2(n_74), .B(n_75), .C(n_78), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_237), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_241), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_250), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_249), .B(n_242), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_260), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_258), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_247), .B(n_235), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_262), .B(n_259), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_261), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_263), .Y(n_268) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_264), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_267), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_271), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_270), .B(n_268), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_272), .Y(n_274) );
NOR2x1p5_ASAP7_75t_L g275 ( .A(n_274), .B(n_273), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_275), .B(n_266), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_276), .B(n_266), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_277), .B(n_266), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_278), .A2(n_257), .B(n_255), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g280 ( .A1(n_279), .A2(n_256), .B1(n_246), .B2(n_251), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g281 ( .A(n_280), .B(n_252), .C(n_253), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_281), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_282), .A2(n_254), .B(n_231), .Y(n_283) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_283), .A2(n_248), .B(n_265), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_284), .B(n_86), .Y(n_285) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_285), .A2(n_87), .B(n_88), .Y(n_286) );
endmodule