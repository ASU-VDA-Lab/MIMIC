module fake_jpeg_16282_n_25 (n_3, n_2, n_1, n_0, n_4, n_5, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_12),
.B1(n_2),
.B2(n_7),
.Y(n_15)
);

OAI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_10),
.C(n_15),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_18),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_10),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_22),
.B(n_10),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_3),
.B(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_25)
);


endmodule