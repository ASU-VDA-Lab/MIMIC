module real_jpeg_29862_n_18 (n_17, n_8, n_0, n_2, n_10, n_338, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_338;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_0),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_0),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_0),
.A2(n_26),
.B1(n_56),
.B2(n_57),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_3),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_5),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_28),
.B(n_32),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_5),
.B(n_30),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_56),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_56),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_68),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_132),
.B1(n_200),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_31),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_6),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_106),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_106),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_9),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_97),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_10),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_100),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_286)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_92),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_92),
.Y(n_220)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_66)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_90),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_90),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_90),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_16),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_16),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_278)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_17),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_25),
.A2(n_34),
.B(n_104),
.C(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_27),
.A2(n_30),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_27),
.A2(n_30),
.B1(n_142),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_27),
.A2(n_30),
.B1(n_161),
.B2(n_258),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_31),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_63),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_31),
.A2(n_57),
.A3(n_217),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_32),
.B(n_104),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_38),
.A2(n_39),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_59),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_40),
.B(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_286),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_46),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_46),
.A2(n_59),
.B1(n_312),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_58),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_54),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_54),
.B1(n_130),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_47),
.A2(n_54),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_47),
.A2(n_54),
.B1(n_175),
.B2(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_47),
.B(n_104),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_47),
.A2(n_54),
.B1(n_96),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_47),
.A2(n_54),
.B1(n_58),
.B2(n_267),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_48),
.A2(n_51),
.A3(n_56),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_49),
.B(n_50),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_50),
.B(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_56),
.B(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_59),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_68),
.B1(n_89),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_61),
.A2(n_68),
.B1(n_145),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_61),
.A2(n_68),
.B1(n_163),
.B2(n_260),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_66),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_66),
.B1(n_88),
.B2(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_62),
.A2(n_66),
.B1(n_91),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_62),
.A2(n_66),
.B1(n_121),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_62),
.A2(n_66),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_69),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_73),
.A2(n_75),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_73),
.A2(n_75),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_327),
.B(n_333),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_303),
.A3(n_322),
.B1(n_325),
.B2(n_326),
.C(n_337),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_254),
.A3(n_292),
.B1(n_297),
.B2(n_302),
.C(n_338),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_147),
.C(n_165),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_125),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_83),
.B(n_125),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_107),
.C(n_117),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_84),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_102),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_94),
.C(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_98),
.A2(n_101),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_98),
.A2(n_101),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_115),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_107),
.A2(n_117),
.B1(n_118),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_107),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_110),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_111),
.A2(n_114),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g270 ( 
.A(n_114),
.Y(n_270)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_119),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_122),
.B(n_124),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_123),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_136),
.C(n_137),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_134),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_132),
.A2(n_134),
.B1(n_194),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_132),
.A2(n_134),
.B1(n_189),
.B2(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_132),
.A2(n_154),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_148),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_149),
.B(n_150),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_152),
.B(n_157),
.C(n_164),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_153),
.B(n_155),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_156),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_248),
.B(n_253),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_234),
.B(n_247),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_210),
.B(n_233),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_190),
.B(n_209),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_170),
.B(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_188),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_197),
.B(n_208),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_207),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_223),
.B1(n_231),
.B2(n_232),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_222),
.C(n_232),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_229),
.Y(n_242)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.C(n_271),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_262),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_256),
.Y(n_335)
);

FAx1_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.CI(n_261),
.CON(n_256),
.SN(n_256)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_258),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_268),
.B2(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_269),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_284),
.B(n_287),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_290),
.B2(n_291),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_281),
.C(n_291),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B(n_280),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_279),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_305),
.C(n_314),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_280),
.B(n_305),
.CI(n_314),
.CON(n_324),
.SN(n_324)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_315),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_313),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_307),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_320),
.C(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule