module fake_jpeg_7773_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_40),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_23),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_28),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_60),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_26),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_62),
.B1(n_66),
.B2(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_22),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_24),
.B1(n_33),
.B2(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_41),
.B1(n_43),
.B2(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_78),
.B1(n_48),
.B2(n_47),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_51),
.B(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_74),
.A2(n_84),
.B1(n_86),
.B2(n_96),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_40),
.A3(n_31),
.B1(n_43),
.B2(n_38),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_95),
.A3(n_82),
.B1(n_54),
.B2(n_91),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_62),
.B1(n_53),
.B2(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_38),
.CI(n_37),
.CON(n_91),
.SN(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_35),
.B1(n_40),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_113),
.B1(n_88),
.B2(n_47),
.Y(n_135)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_106),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_117),
.Y(n_134)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_61),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_65),
.C(n_30),
.Y(n_148)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_115),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_47),
.B1(n_55),
.B2(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_49),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_70),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_94),
.B(n_89),
.C(n_49),
.D(n_65),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_70),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_69),
.B1(n_49),
.B2(n_64),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_122),
.B1(n_115),
.B2(n_110),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_75),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_136),
.B(n_98),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_78),
.B1(n_90),
.B2(n_91),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_135),
.Y(n_154)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_71),
.B(n_84),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_74),
.B1(n_90),
.B2(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_94),
.B1(n_89),
.B2(n_69),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_143),
.B1(n_152),
.B2(n_101),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_103),
.Y(n_168)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_47),
.B1(n_72),
.B2(n_81),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_108),
.C(n_117),
.Y(n_157)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_81),
.B1(n_55),
.B2(n_58),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_77),
.B1(n_52),
.B2(n_50),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_41),
.B1(n_30),
.B2(n_17),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_158),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_160),
.C(n_179),
.Y(n_186)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

OAI22x1_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_121),
.B1(n_125),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_123),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_140),
.C(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_116),
.B(n_107),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_180),
.B(n_25),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_116),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_103),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_25),
.CI(n_38),
.CON(n_206),
.SN(n_206)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_104),
.B1(n_114),
.B2(n_120),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_106),
.B1(n_41),
.B2(n_17),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_38),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_0),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_20),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_150),
.B1(n_131),
.B2(n_137),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_130),
.B1(n_145),
.B2(n_127),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_185),
.B(n_199),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_153),
.B(n_144),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_147),
.C(n_148),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_147),
.C(n_139),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_134),
.C(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_200),
.B1(n_32),
.B2(n_23),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_159),
.A2(n_152),
.B(n_25),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_182),
.B1(n_154),
.B2(n_172),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_141),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_77),
.C(n_52),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_18),
.C(n_21),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_38),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_38),
.C(n_50),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_171),
.B(n_170),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_211),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_161),
.C(n_166),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_164),
.B1(n_169),
.B2(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_218),
.B1(n_219),
.B2(n_223),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_216),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_180),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_235),
.C(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_180),
.B(n_178),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_231),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_169),
.B1(n_177),
.B2(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_173),
.B1(n_141),
.B2(n_23),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_52),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_226),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_27),
.B1(n_23),
.B2(n_32),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_50),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_18),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_208),
.Y(n_245)
);

NOR4xp25_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_12),
.C(n_9),
.D(n_16),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_18),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_184),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_198),
.A2(n_12),
.B(n_16),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_199),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_12),
.C(n_15),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_7),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_240),
.C(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_195),
.C(n_184),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_188),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.C(n_254),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_192),
.C(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.C(n_33),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_192),
.C(n_183),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_233),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_266),
.C(n_269),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_183),
.B1(n_210),
.B2(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_264),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_230),
.CI(n_218),
.CON(n_264),
.SN(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_235),
.B1(n_32),
.B2(n_27),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_33),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_18),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_32),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_27),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_27),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_253),
.B(n_7),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_236),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_33),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_238),
.B(n_246),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_275),
.A2(n_13),
.B(n_10),
.Y(n_301)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_239),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_285),
.B(n_286),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_254),
.CI(n_242),
.CON(n_279),
.SN(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_289),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_249),
.C(n_245),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_271),
.C(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_268),
.B1(n_274),
.B2(n_271),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_276),
.A3(n_279),
.B1(n_284),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_294),
.C(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_266),
.C(n_21),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_275),
.B1(n_276),
.B2(n_279),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_1),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_14),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_2),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_281),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_302),
.B(n_2),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_13),
.B(n_10),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_307),
.B1(n_312),
.B2(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_2),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_310),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_291),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_297),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_300),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_320),
.B(n_292),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_323),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_3),
.B(n_4),
.Y(n_324)
);

AOI321xp33_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_5),
.A3(n_6),
.B1(n_318),
.B2(n_320),
.C(n_322),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_5),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_5),
.Y(n_328)
);

XNOR2x2_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_6),
.Y(n_329)
);


endmodule