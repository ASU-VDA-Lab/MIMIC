module fake_jpeg_19834_n_100 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_12),
.B(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_15),
.B1(n_31),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_18),
.Y(n_61)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_11),
.B1(n_29),
.B2(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_33),
.B1(n_27),
.B2(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_54),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_39),
.B1(n_35),
.B2(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_60),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_24),
.B(n_19),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_65),
.B(n_0),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_54),
.B1(n_51),
.B2(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_0),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_71),
.B(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_3),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_82),
.B(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_84),
.B1(n_68),
.B2(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_80),
.A2(n_68),
.B1(n_66),
.B2(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_89),
.B1(n_81),
.B2(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_58),
.B1(n_62),
.B2(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_83),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.C(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_89),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_7),
.B(n_8),
.Y(n_97)
);

AOI31xp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_9),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_10),
.B(n_72),
.Y(n_100)
);


endmodule