module fake_jpeg_13486_n_76 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_76);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_76;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_25),
.B2(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_14),
.B(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_3),
.Y(n_55)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_4),
.C(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_11),
.B1(n_19),
.B2(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.C(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_55),
.C(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_63),
.Y(n_70)
);

XNOR2x1_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_69),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_62),
.B(n_16),
.Y(n_74)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_15),
.B(n_17),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_18),
.CI(n_24),
.CON(n_76),
.SN(n_76)
);


endmodule