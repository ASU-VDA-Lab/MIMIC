module real_jpeg_25989_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_0),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_5),
.A2(n_20),
.B1(n_26),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_25),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_25),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_6),
.B(n_52),
.C(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_33),
.C(n_47),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_20),
.C(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_6),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_106),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_104),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_90),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_90),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_68),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_42),
.B(n_65),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_16),
.A2(n_17),
.B1(n_70),
.B2(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_31),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_18),
.A2(n_31),
.B1(n_93),
.B2(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_19),
.A2(n_29),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_20),
.B(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_31),
.A2(n_73),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_31),
.Y(n_93)
);

AOI211xp5_ASAP7_75t_L g113 ( 
.A1(n_31),
.A2(n_55),
.B(n_65),
.C(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_31),
.A2(n_44),
.B1(n_67),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_31),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_31),
.A2(n_93),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_31),
.A2(n_93),
.B1(n_147),
.B2(n_148),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_31),
.A2(n_44),
.B(n_114),
.C(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_31),
.A2(n_93),
.B1(n_135),
.B2(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_33),
.B(n_149),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_37),
.A2(n_40),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_96),
.B(n_103),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_55),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_44),
.B(n_97),
.C(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_44),
.A2(n_67),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_46),
.Y(n_155)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_52),
.B(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_66),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_78),
.B1(n_88),
.B2(n_89),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_71),
.B1(n_96),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.C(n_95),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_91),
.B(n_92),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_132),
.C(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_93),
.B(n_98),
.C(n_154),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_95),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_98),
.B1(n_125),
.B2(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_97),
.A2(n_98),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_97),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_97),
.A2(n_98),
.B1(n_136),
.B2(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_98),
.B(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_128),
.B(n_182),
.C(n_186),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_118),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_117),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_113),
.C(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_121),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_181),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_142),
.B(n_180),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_139),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_131),
.B(n_139),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_174),
.B(n_179),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_168),
.B(n_173),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_156),
.B(n_167),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.Y(n_186)
);


endmodule