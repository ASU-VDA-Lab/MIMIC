module fake_ibex_1453_n_1159 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1159);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1159;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1148;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1018;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1138;
wire n_727;
wire n_1134;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_280;
wire n_340;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_1109;
wire n_210;
wire n_348;
wire n_965;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_497;
wire n_287;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_1057;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_234;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_1092;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_209;
wire n_229;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_940;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_1150;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_890;
wire n_816;
wire n_874;
wire n_912;
wire n_1058;
wire n_1105;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_76),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_23),
.B(n_57),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_80),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_130),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_30),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_119),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_29),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_165),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_111),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_43),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_126),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_185),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_70),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_208),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_39),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_161),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_143),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_34),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_34),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_69),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_188),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_98),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_66),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_191),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_181),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_147),
.B(n_40),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_136),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_135),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_41),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_68),
.Y(n_273)
);

BUFx2_ASAP7_75t_SL g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_113),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_77),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_121),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_138),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_102),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_116),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_129),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_24),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_171),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_81),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_115),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_38),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_174),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_179),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_200),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_132),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_3),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_131),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_55),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_112),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_87),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_122),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_108),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_199),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_159),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_139),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_158),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_85),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_33),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_95),
.B(n_196),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_11),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_14),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_38),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_93),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_86),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_190),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_197),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_169),
.Y(n_321)
);

BUFx2_ASAP7_75t_SL g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_83),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_92),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_182),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_203),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_37),
.B(n_48),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_29),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_180),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_10),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_173),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_177),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_48),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_15),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_193),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_110),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_28),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_60),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_155),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_120),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_192),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_25),
.B(n_35),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_142),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_44),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_101),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_8),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_84),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_60),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_107),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_117),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_178),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_118),
.B(n_114),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_72),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_2),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_176),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_128),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_163),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_18),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_16),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_194),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_21),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_96),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_39),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_187),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_41),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_146),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_52),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_256),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_231),
.Y(n_374)
);

BUFx8_ASAP7_75t_SL g375 ( 
.A(n_218),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_269),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_243),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_211),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_316),
.B(n_0),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_63),
.Y(n_383)
);

BUFx12f_ASAP7_75t_L g384 ( 
.A(n_223),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_210),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_210),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_218),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_210),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_222),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_290),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_223),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_290),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_222),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_225),
.A2(n_65),
.B(n_64),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_271),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_253),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_222),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_271),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_291),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_230),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_299),
.B(n_1),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_258),
.B(n_3),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_292),
.Y(n_409)
);

BUFx8_ASAP7_75t_SL g410 ( 
.A(n_286),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_230),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_222),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_230),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_230),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_230),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_289),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_230),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_318),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_289),
.Y(n_422)
);

AOI22x1_ASAP7_75t_SL g423 ( 
.A1(n_306),
.A2(n_320),
.B1(n_331),
.B2(n_309),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_223),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_230),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_289),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_289),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_300),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_300),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_211),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_209),
.B(n_212),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_247),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_302),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_300),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_228),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_300),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_227),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_262),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_225),
.A2(n_99),
.B(n_205),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_302),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_262),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_278),
.A2(n_97),
.B(n_204),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_224),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_258),
.B(n_12),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_213),
.B(n_12),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_343),
.B(n_325),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_302),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_325),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_232),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_236),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_362),
.B(n_13),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_238),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_248),
.Y(n_454)
);

OAI22x1_ASAP7_75t_SL g455 ( 
.A1(n_309),
.A2(n_331),
.B1(n_333),
.B2(n_320),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_224),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_259),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_254),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_333),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_362),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_281),
.Y(n_461)
);

INVx6_ASAP7_75t_L g462 ( 
.A(n_302),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_282),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_302),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_343),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_266),
.B(n_311),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_314),
.B(n_17),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_302),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_282),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_295),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_255),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_381),
.B(n_373),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_261),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_406),
.B(n_360),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_394),
.B(n_301),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_405),
.B(n_272),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_374),
.B(n_275),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_400),
.A2(n_339),
.B1(n_335),
.B2(n_329),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_406),
.B(n_360),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_376),
.B(n_297),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_217),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

NOR2x1_ASAP7_75t_L g488 ( 
.A(n_377),
.B(n_219),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_L g490 ( 
.A(n_383),
.B(n_357),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_400),
.B(n_317),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_452),
.B(n_233),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_330),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_402),
.B(n_332),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_237),
.Y(n_497)
);

NOR2x1p5_ASAP7_75t_L g498 ( 
.A(n_384),
.B(n_351),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_436),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_SL g500 ( 
.A(n_408),
.B(n_339),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_SL g501 ( 
.A(n_408),
.B(n_215),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_L g502 ( 
.A1(n_402),
.A2(n_359),
.B1(n_363),
.B2(n_353),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_438),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_375),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_445),
.B(n_220),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_383),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_461),
.B(n_250),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_463),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_404),
.B(n_337),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_439),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_380),
.B(n_341),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_382),
.B(n_344),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_461),
.B(n_252),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_439),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_379),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_465),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_458),
.B(n_368),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_439),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_442),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_466),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_214),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_268),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_472),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_431),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_442),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_419),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_450),
.B(n_270),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_280),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_461),
.B(n_283),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_453),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_457),
.B(n_288),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_461),
.B(n_296),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_383),
.B(n_221),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_388),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_460),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

INVxp33_ASAP7_75t_L g560 ( 
.A(n_386),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_409),
.B(n_308),
.Y(n_561)
);

INVxp67_ASAP7_75t_R g562 ( 
.A(n_455),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_393),
.A2(n_366),
.B1(n_364),
.B2(n_235),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_411),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_445),
.B(n_284),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_399),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_413),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g569 ( 
.A1(n_443),
.A2(n_321),
.B(n_319),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_403),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_415),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_416),
.B(n_324),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_416),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_449),
.B(n_226),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_425),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_425),
.B(n_427),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_427),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_434),
.B(n_345),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_441),
.B(n_348),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_448),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_420),
.B(n_350),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_388),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_410),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_469),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_414),
.A2(n_313),
.B1(n_349),
.B2(n_342),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_410),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_421),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_397),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_385),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_421),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_421),
.B(n_234),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_558),
.A2(n_432),
.B1(n_459),
.B2(n_446),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_594),
.Y(n_601)
);

AO221x1_ASAP7_75t_L g602 ( 
.A1(n_483),
.A2(n_423),
.B1(n_241),
.B2(n_245),
.C(n_249),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_597),
.Y(n_603)
);

NOR2xp67_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_506),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_560),
.B(n_274),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_473),
.A2(n_251),
.B1(n_293),
.B2(n_265),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_354),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_560),
.A2(n_371),
.B1(n_328),
.B2(n_347),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_529),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_239),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_546),
.B(n_240),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_523),
.B(n_242),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_526),
.B(n_244),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_597),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_495),
.B(n_358),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_597),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_246),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_522),
.B(n_322),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_539),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_504),
.B(n_257),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_492),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_555),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_535),
.B(n_369),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_478),
.B(n_486),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_593),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_497),
.B(n_229),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_512),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_590),
.B(n_216),
.C(n_263),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_496),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_513),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_522),
.B(n_224),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_599),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_567),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_536),
.B(n_488),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

AO221x1_ASAP7_75t_L g642 ( 
.A1(n_502),
.A2(n_444),
.B1(n_456),
.B2(n_426),
.C(n_437),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_503),
.A2(n_352),
.B1(n_267),
.B2(n_273),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_474),
.A2(n_355),
.B1(n_276),
.B2(n_277),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_481),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_490),
.B(n_440),
.C(n_397),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_R g647 ( 
.A(n_552),
.B(n_500),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_548),
.B(n_279),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_485),
.B(n_287),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_520),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_519),
.B(n_264),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_542),
.B(n_294),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_543),
.B(n_298),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_480),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_482),
.B(n_305),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_285),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_509),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_531),
.B(n_307),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_493),
.B(n_310),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_595),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_561),
.B(n_323),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_547),
.B(n_327),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_598),
.B(n_338),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_499),
.B(n_340),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_537),
.B(n_346),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_477),
.B(n_356),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_490),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_505),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_576),
.B(n_361),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_584),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_551),
.A2(n_444),
.B1(n_456),
.B2(n_437),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_484),
.B(n_367),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_564),
.B(n_19),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_498),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_525),
.B(n_312),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_508),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_500),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_574),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_525),
.B(n_534),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_541),
.B(n_20),
.Y(n_685)
);

AO221x1_ASAP7_75t_L g686 ( 
.A1(n_494),
.A2(n_456),
.B1(n_437),
.B2(n_378),
.C(n_430),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_573),
.B(n_565),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_501),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_501),
.A2(n_456),
.B1(n_417),
.B2(n_412),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_574),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_534),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_585),
.B(n_21),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_568),
.B(n_417),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_516),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_507),
.A2(n_417),
.B1(n_430),
.B2(n_429),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_571),
.B(n_378),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_581),
.B(n_387),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_572),
.B(n_389),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_596),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_575),
.B(n_577),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_646),
.A2(n_579),
.B(n_569),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_628),
.A2(n_582),
.B(n_592),
.C(n_589),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_608),
.B(n_588),
.C(n_524),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_682),
.A2(n_583),
.B1(n_592),
.B2(n_575),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_691),
.B(n_591),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_628),
.B(n_580),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_659),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_601),
.B(n_511),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_664),
.A2(n_550),
.B(n_545),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_659),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_639),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_625),
.B(n_591),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_605),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_607),
.A2(n_586),
.B(n_587),
.C(n_476),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_675),
.B(n_627),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_699),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_625),
.A2(n_491),
.B1(n_489),
.B2(n_479),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_653),
.B(n_487),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_672),
.A2(n_527),
.B1(n_563),
.B2(n_557),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_637),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_623),
.A2(n_634),
.B(n_645),
.C(n_635),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_623),
.B(n_22),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_658),
.B(n_616),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_658),
.B(n_22),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_687),
.A2(n_700),
.B(n_672),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_616),
.B(n_23),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_647),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_656),
.A2(n_690),
.B(n_683),
.Y(n_729)
);

OAI321xp33_ASAP7_75t_L g730 ( 
.A1(n_608),
.A2(n_435),
.A3(n_401),
.B1(n_396),
.B2(n_390),
.C(n_389),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_688),
.A2(n_540),
.B1(n_517),
.B2(n_556),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_633),
.A2(n_563),
.B1(n_517),
.B2(n_556),
.Y(n_732)
);

CKINVDCx8_ASAP7_75t_R g733 ( 
.A(n_670),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_651),
.A2(n_532),
.B(n_554),
.C(n_553),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_685),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_641),
.B(n_25),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_678),
.B(n_26),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_640),
.B(n_26),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_632),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_619),
.B(n_27),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_600),
.A2(n_532),
.B1(n_549),
.B2(n_544),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_631),
.B(n_31),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_610),
.B(n_31),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_633),
.A2(n_518),
.B(n_527),
.C(n_528),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_604),
.B(n_533),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_612),
.A2(n_618),
.B(n_614),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_677),
.A2(n_538),
.B(n_35),
.C(n_36),
.Y(n_748)
);

BUFx4f_ASAP7_75t_L g749 ( 
.A(n_692),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_609),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_689),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_652),
.B(n_32),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_660),
.B(n_661),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_679),
.B(n_42),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_671),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_657),
.B(n_636),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_630),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_666),
.B(n_46),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_650),
.B(n_47),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_654),
.B(n_49),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_684),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_R g762 ( 
.A(n_655),
.B(n_49),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_603),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_695),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_662),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_648),
.B(n_644),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_663),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_50),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_615),
.A2(n_617),
.B(n_697),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_667),
.B(n_669),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_621),
.A2(n_626),
.B(n_622),
.C(n_629),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_668),
.B(n_51),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_642),
.A2(n_429),
.B1(n_428),
.B2(n_426),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_697),
.A2(n_401),
.B(n_428),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_624),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_674),
.A2(n_422),
.B(n_396),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_680),
.B(n_56),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_665),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_638),
.A2(n_422),
.B1(n_396),
.B2(n_59),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_611),
.A2(n_422),
.B(n_124),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_686),
.B(n_57),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_676),
.B(n_61),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_693),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_602),
.B(n_202),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_724),
.B(n_696),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_775),
.A2(n_698),
.A3(n_681),
.B(n_694),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_712),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_711),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_716),
.B(n_673),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_738),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_757),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_705),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_710),
.B(n_737),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_710),
.B(n_740),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_706),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_705),
.Y(n_797)
);

AOI21xp33_ASAP7_75t_L g798 ( 
.A1(n_722),
.A2(n_753),
.B(n_714),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_756),
.A2(n_88),
.B(n_89),
.C(n_90),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_707),
.B(n_91),
.Y(n_800)
);

AO31x2_ASAP7_75t_L g801 ( 
.A1(n_734),
.A2(n_100),
.A3(n_106),
.B(n_109),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_762),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_705),
.Y(n_803)
);

BUFx4_ASAP7_75t_SL g804 ( 
.A(n_728),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_723),
.B(n_140),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_735),
.B(n_141),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_726),
.A2(n_144),
.B(n_148),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_713),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_741),
.B(n_766),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_702),
.A2(n_157),
.B(n_160),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_703),
.A2(n_166),
.B1(n_167),
.B2(n_170),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_729),
.A2(n_172),
.B(n_175),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_736),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_765),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_771),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_719),
.B(n_721),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_776),
.A2(n_743),
.B(n_744),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_749),
.B(n_733),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_758),
.B(n_760),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_771),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_SL g822 ( 
.A1(n_715),
.A2(n_748),
.B(n_745),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_771),
.Y(n_823)
);

NAND2x1_ASAP7_75t_L g824 ( 
.A(n_717),
.B(n_767),
.Y(n_824)
);

AO21x2_ASAP7_75t_L g825 ( 
.A1(n_730),
.A2(n_769),
.B(n_777),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_708),
.B(n_727),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_765),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_725),
.A2(n_755),
.B(n_759),
.C(n_773),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_708),
.B(n_768),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_739),
.B(n_718),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_717),
.B(n_779),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_772),
.A2(n_709),
.B(n_763),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_746),
.Y(n_833)
);

OAI21x1_ASAP7_75t_SL g834 ( 
.A1(n_774),
.A2(n_778),
.B(n_767),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_754),
.B(n_761),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_784),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_751),
.B(n_704),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_764),
.A2(n_785),
.B1(n_732),
.B2(n_783),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_720),
.A2(n_742),
.B(n_781),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_750),
.A2(n_770),
.B1(n_780),
.B2(n_731),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_705),
.B(n_649),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_706),
.A2(n_672),
.B1(n_716),
.B2(n_724),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_724),
.B(n_716),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_724),
.B(n_716),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_706),
.A2(n_724),
.B1(n_716),
.B2(n_672),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_710),
.B(n_649),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_710),
.B(n_560),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_724),
.A2(n_747),
.B(n_716),
.C(n_628),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_724),
.B(n_716),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_737),
.B(n_494),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_710),
.B(n_560),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_705),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_724),
.B(n_716),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_724),
.B(n_716),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_701),
.A2(n_646),
.B(n_726),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_560),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_712),
.Y(n_857)
);

AO31x2_ASAP7_75t_L g858 ( 
.A1(n_775),
.A2(n_701),
.A3(n_782),
.B(n_595),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_710),
.B(n_649),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_724),
.A2(n_747),
.B(n_716),
.C(n_628),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_724),
.B(n_716),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_711),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_710),
.B(n_649),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_724),
.B(n_716),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_724),
.B(n_716),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_737),
.B(n_494),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_712),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_724),
.B(n_716),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_705),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_712),
.B(n_757),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_701),
.A2(n_646),
.B(n_726),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_712),
.Y(n_872)
);

AOI221xp5_ASAP7_75t_SL g873 ( 
.A1(n_745),
.A2(n_748),
.B1(n_716),
.B2(n_724),
.C(n_727),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_710),
.B(n_649),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_724),
.B(n_716),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_724),
.B(n_716),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_724),
.B(n_716),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_701),
.A2(n_490),
.B(n_551),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_724),
.B(n_716),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_710),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_710),
.B(n_560),
.Y(n_881)
);

BUFx10_ASAP7_75t_L g882 ( 
.A(n_705),
.Y(n_882)
);

AND3x4_ASAP7_75t_L g883 ( 
.A(n_703),
.B(n_604),
.C(n_562),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_724),
.B(n_716),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_705),
.Y(n_885)
);

AO31x2_ASAP7_75t_L g886 ( 
.A1(n_775),
.A2(n_701),
.A3(n_782),
.B(n_595),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_724),
.B(n_716),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_706),
.A2(n_724),
.B1(n_716),
.B2(n_672),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_712),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_701),
.A2(n_646),
.B(n_726),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_710),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_859),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_848),
.A2(n_860),
.B(n_842),
.Y(n_893)
);

INVx3_ASAP7_75t_SL g894 ( 
.A(n_852),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_815),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_815),
.B(n_827),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_792),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_842),
.Y(n_898)
);

AO21x2_ASAP7_75t_L g899 ( 
.A1(n_871),
.A2(n_890),
.B(n_834),
.Y(n_899)
);

CKINVDCx11_ASAP7_75t_R g900 ( 
.A(n_869),
.Y(n_900)
);

BUFx2_ASAP7_75t_SL g901 ( 
.A(n_793),
.Y(n_901)
);

BUFx2_ASAP7_75t_SL g902 ( 
.A(n_793),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_838),
.B(n_811),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_880),
.B(n_863),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_843),
.B(n_844),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_827),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_841),
.B(n_885),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_870),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_841),
.B(n_833),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_849),
.B(n_853),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_870),
.Y(n_912)
);

CKINVDCx6p67_ASAP7_75t_R g913 ( 
.A(n_841),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_882),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_847),
.B(n_851),
.Y(n_915)
);

CKINVDCx11_ASAP7_75t_R g916 ( 
.A(n_882),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_788),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_873),
.B(n_828),
.C(n_810),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_878),
.A2(n_888),
.B(n_845),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_856),
.Y(n_920)
);

CKINVDCx6p67_ASAP7_75t_R g921 ( 
.A(n_797),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_870),
.B(n_854),
.Y(n_922)
);

BUFx4_ASAP7_75t_SL g923 ( 
.A(n_816),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_861),
.B(n_864),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_881),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_839),
.A2(n_822),
.B(n_825),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_865),
.B(n_868),
.Y(n_927)
);

NOR2x1_ASAP7_75t_R g928 ( 
.A(n_802),
.B(n_821),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_891),
.Y(n_929)
);

NOR2x1_ASAP7_75t_SL g930 ( 
.A(n_875),
.B(n_876),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_836),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_804),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_857),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_825),
.A2(n_832),
.B(n_807),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_798),
.A2(n_794),
.B1(n_809),
.B2(n_837),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_877),
.B(n_879),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_831),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_884),
.B(n_887),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_823),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_867),
.B(n_872),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_796),
.A2(n_813),
.B(n_811),
.Y(n_941)
);

NOR2x1_ASAP7_75t_R g942 ( 
.A(n_803),
.B(n_819),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_889),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_830),
.A2(n_791),
.B1(n_817),
.B2(n_805),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_824),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_826),
.A2(n_786),
.B(n_829),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_840),
.A2(n_806),
.B(n_796),
.Y(n_947)
);

AO31x2_ASAP7_75t_L g948 ( 
.A1(n_840),
.A2(n_799),
.A3(n_886),
.B(n_858),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_791),
.A2(n_814),
.B(n_818),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_795),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_820),
.A2(n_812),
.B(n_790),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_850),
.B(n_866),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_835),
.B(n_808),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_846),
.B(n_874),
.Y(n_954)
);

XNOR2xp5_ASAP7_75t_L g955 ( 
.A(n_883),
.B(n_800),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_787),
.A2(n_858),
.B(n_886),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_787),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_787),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_801),
.A2(n_862),
.B(n_855),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_815),
.B(n_827),
.Y(n_960)
);

BUFx8_ASAP7_75t_L g961 ( 
.A(n_869),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_880),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_841),
.B(n_869),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_870),
.B(n_843),
.Y(n_964)
);

CKINVDCx6p67_ASAP7_75t_R g965 ( 
.A(n_852),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_848),
.A2(n_860),
.B(n_842),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_804),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_815),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_927),
.B(n_936),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_940),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_905),
.B(n_911),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_940),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_931),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_912),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_927),
.B(n_930),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_917),
.Y(n_976)
);

AO21x1_ASAP7_75t_SL g977 ( 
.A1(n_893),
.A2(n_966),
.B(n_919),
.Y(n_977)
);

CKINVDCx11_ASAP7_75t_R g978 ( 
.A(n_894),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_931),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_908),
.B(n_947),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_933),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_905),
.B(n_911),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_943),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_899),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_899),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_896),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_SL g987 ( 
.A1(n_944),
.A2(n_922),
.B1(n_964),
.B2(n_901),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_924),
.B(n_938),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_932),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_924),
.B(n_938),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_SL g991 ( 
.A1(n_898),
.A2(n_903),
.B(n_893),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_957),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_937),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_950),
.B(n_935),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_958),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_961),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_897),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_952),
.A2(n_964),
.B1(n_935),
.B2(n_925),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_SL g999 ( 
.A1(n_902),
.A2(n_929),
.B1(n_898),
.B2(n_952),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_923),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_953),
.A2(n_920),
.B1(n_941),
.B2(n_915),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_959),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_895),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_953),
.A2(n_946),
.B1(n_951),
.B2(n_949),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_909),
.Y(n_1005)
);

OAI22xp33_ASAP7_75t_SL g1006 ( 
.A1(n_962),
.A2(n_968),
.B1(n_906),
.B2(n_895),
.Y(n_1006)
);

BUFx2_ASAP7_75t_R g1007 ( 
.A(n_967),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_999),
.B(n_892),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_977),
.B(n_956),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_977),
.B(n_926),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_1005),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_970),
.B(n_918),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_972),
.B(n_918),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_992),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_992),
.B(n_926),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_995),
.B(n_948),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_995),
.B(n_948),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_1003),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_973),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_994),
.B(n_906),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_991),
.B(n_948),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_991),
.B(n_934),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_979),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_976),
.Y(n_1025)
);

INVx3_ASAP7_75t_SL g1026 ( 
.A(n_993),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_996),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_1005),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_975),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_981),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_1005),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_969),
.B(n_960),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1001),
.A2(n_962),
.B1(n_913),
.B2(n_910),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1014),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1014),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1025),
.B(n_982),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_L g1038 ( 
.A(n_1017),
.B(n_986),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1015),
.B(n_1016),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1021),
.B(n_969),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1025),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1009),
.B(n_980),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1017),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_1033),
.A2(n_987),
.B1(n_982),
.B2(n_988),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1021),
.B(n_1004),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1019),
.B(n_984),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1015),
.B(n_985),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1015),
.B(n_985),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1020),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1016),
.B(n_1002),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_1017),
.B(n_974),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1020),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1033),
.A2(n_988),
.B1(n_971),
.B2(n_998),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1039),
.B(n_1019),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1039),
.B(n_1010),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1050),
.B(n_1010),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1050),
.B(n_1047),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1049),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1035),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_1043),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1035),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1052),
.Y(n_1062)
);

NAND4xp25_ASAP7_75t_L g1063 ( 
.A(n_1044),
.B(n_990),
.C(n_1008),
.D(n_1010),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1047),
.B(n_1009),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1036),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1042),
.B(n_1009),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1036),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_L g1068 ( 
.A(n_1051),
.B(n_1000),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1037),
.B(n_1024),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1034),
.B(n_1024),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1034),
.B(n_1030),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1041),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1048),
.B(n_1016),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_1043),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1054),
.Y(n_1075)
);

INVxp33_ASAP7_75t_L g1076 ( 
.A(n_1054),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1058),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1062),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1059),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1057),
.B(n_1042),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1070),
.B(n_1045),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1059),
.Y(n_1082)
);

NAND2x1_ASAP7_75t_L g1083 ( 
.A(n_1066),
.B(n_1051),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1071),
.B(n_1073),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1061),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1073),
.B(n_1018),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1060),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1057),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1069),
.B(n_1040),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1077),
.B(n_1063),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1075),
.B(n_1055),
.Y(n_1092)
);

AOI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_1076),
.A2(n_1026),
.B(n_894),
.C(n_1000),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1079),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1082),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1088),
.B(n_1055),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1085),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1080),
.B(n_1064),
.Y(n_1098)
);

AOI21xp33_ASAP7_75t_SL g1099 ( 
.A1(n_1074),
.A2(n_1026),
.B(n_996),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1084),
.B(n_1064),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1078),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1084),
.B(n_1056),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1081),
.A2(n_1053),
.B1(n_1056),
.B2(n_1067),
.C(n_1072),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1074),
.A2(n_1038),
.B(n_975),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1090),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1074),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1091),
.A2(n_1089),
.B1(n_1066),
.B2(n_1083),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_SL g1108 ( 
.A(n_1099),
.B(n_1087),
.C(n_1027),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1091),
.A2(n_1089),
.B1(n_1086),
.B2(n_1042),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1093),
.A2(n_1089),
.B(n_1006),
.Y(n_1110)
);

AOI222xp33_ASAP7_75t_L g1111 ( 
.A1(n_1103),
.A2(n_1086),
.B1(n_1022),
.B2(n_1023),
.C1(n_1065),
.C2(n_978),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1094),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1104),
.A2(n_1006),
.B(n_1028),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1106),
.A2(n_1026),
.B1(n_1017),
.B2(n_1040),
.Y(n_1114)
);

OAI32xp33_ASAP7_75t_L g1115 ( 
.A1(n_1106),
.A2(n_1029),
.A3(n_1045),
.B1(n_1031),
.B2(n_1011),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1108),
.A2(n_1101),
.B(n_1097),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1107),
.B(n_1105),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1111),
.B(n_1100),
.Y(n_1118)
);

AOI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1114),
.A2(n_928),
.B(n_942),
.Y(n_1119)
);

NAND4xp25_ASAP7_75t_L g1120 ( 
.A(n_1110),
.B(n_954),
.C(n_993),
.D(n_1032),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1112),
.Y(n_1121)
);

OAI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_1109),
.A2(n_1102),
.B(n_1100),
.Y(n_1122)
);

AOI221x1_ASAP7_75t_L g1123 ( 
.A1(n_1113),
.A2(n_1095),
.B1(n_1092),
.B2(n_983),
.C(n_997),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_1115),
.A2(n_1102),
.B1(n_963),
.B2(n_907),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1121),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1116),
.B(n_1098),
.Y(n_1126)
);

AOI32xp33_ASAP7_75t_L g1127 ( 
.A1(n_1118),
.A2(n_1098),
.A3(n_1096),
.B1(n_1029),
.B2(n_1022),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1120),
.A2(n_1117),
.B1(n_1122),
.B2(n_1124),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1123),
.B(n_1096),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1119),
.B(n_961),
.C(n_900),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_SL g1131 ( 
.A(n_1118),
.B(n_1007),
.C(n_989),
.D(n_1032),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1121),
.B(n_1046),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_L g1133 ( 
.A(n_1131),
.B(n_916),
.C(n_993),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_L g1134 ( 
.A(n_1130),
.B(n_904),
.C(n_954),
.Y(n_1134)
);

NOR3x1_ASAP7_75t_L g1135 ( 
.A(n_1126),
.B(n_989),
.C(n_965),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1125),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_L g1137 ( 
.A(n_1129),
.B(n_907),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1128),
.B(n_914),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1132),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1127),
.B(n_1061),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1138),
.B(n_907),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1136),
.B(n_963),
.C(n_910),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1137),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1133),
.B(n_963),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1140),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_1134),
.B(n_939),
.C(n_945),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1135),
.Y(n_1148)
);

INVxp33_ASAP7_75t_SL g1149 ( 
.A(n_1142),
.Y(n_1149)
);

AND2x2_ASAP7_75t_SL g1150 ( 
.A(n_1147),
.B(n_1146),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1149),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1151),
.B(n_1150),
.Y(n_1152)
);

XNOR2xp5_ASAP7_75t_L g1153 ( 
.A(n_1152),
.B(n_1148),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1153),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1154),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1155),
.B(n_1148),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1156),
.B(n_1141),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_1157),
.A2(n_1144),
.B1(n_1143),
.B2(n_955),
.C(n_921),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1158),
.A2(n_910),
.B(n_923),
.Y(n_1159)
);


endmodule