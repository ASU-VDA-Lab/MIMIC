module fake_jpeg_747_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_7),
.B(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_87),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_14),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_62),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_81),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_93),
.B1(n_97),
.B2(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_1),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_90),
.Y(n_129)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_96),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_95),
.Y(n_142)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_6),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_40),
.B1(n_32),
.B2(n_37),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_119),
.B1(n_121),
.B2(n_86),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_28),
.B1(n_40),
.B2(n_47),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_47),
.B1(n_45),
.B2(n_8),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_47),
.C(n_7),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_110),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_62),
.B(n_10),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_53),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_72),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_89),
.Y(n_161)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_148),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx5_ASAP7_75t_SL g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_97),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_164),
.Y(n_188)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_173),
.B1(n_178),
.B2(n_131),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_63),
.B1(n_88),
.B2(n_95),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_124),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_174),
.Y(n_197)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_144),
.B1(n_119),
.B2(n_120),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

BUFx6f_ASAP7_75t_SL g189 ( 
.A(n_170),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_100),
.A2(n_109),
.B1(n_142),
.B2(n_126),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_104),
.A2(n_100),
.B1(n_113),
.B2(n_135),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_123),
.B1(n_126),
.B2(n_143),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_110),
.A2(n_136),
.B(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_106),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_176),
.Y(n_195)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_115),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_143),
.B1(n_102),
.B2(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_102),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_115),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_150),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_152),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_136),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_179),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_163),
.B1(n_154),
.B2(n_158),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_111),
.B1(n_103),
.B2(n_112),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_174),
.B1(n_160),
.B2(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_205),
.B1(n_173),
.B2(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_117),
.B1(n_125),
.B2(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_164),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_218),
.C(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_216),
.B1(n_224),
.B2(n_190),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_156),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_219),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_153),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_148),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_166),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_176),
.B1(n_170),
.B2(n_132),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_205),
.B1(n_191),
.B2(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_108),
.B1(n_112),
.B2(n_149),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_159),
.B1(n_167),
.B2(n_103),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_201),
.B1(n_186),
.B2(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_238),
.C(n_218),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_190),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_241),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_237),
.B(n_227),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_188),
.B1(n_186),
.B2(n_192),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_183),
.C(n_194),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_194),
.B1(n_183),
.B2(n_196),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_192),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_259),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_216),
.B1(n_222),
.B2(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_228),
.B1(n_220),
.B2(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_213),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_218),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_260),
.Y(n_262)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_218),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_251),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_231),
.B1(n_237),
.B2(n_240),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_272),
.B1(n_248),
.B2(n_255),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_246),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_212),
.B1(n_250),
.B2(n_254),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_274),
.A2(n_268),
.B(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_252),
.C(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_273),
.C(n_262),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_270),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_260),
.B1(n_212),
.B2(n_217),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_235),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_277),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_267),
.B(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

OAI322xp33_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_243),
.A3(n_245),
.B1(n_267),
.B2(n_235),
.C1(n_217),
.C2(n_225),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_208),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_296),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_276),
.B1(n_275),
.B2(n_282),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_299),
.B1(n_292),
.B2(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_284),
.C(n_275),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_245),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_239),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_232),
.B(n_239),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_267),
.B1(n_291),
.B2(n_296),
.Y(n_303)
);

INVx11_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_226),
.A3(n_139),
.B1(n_184),
.B2(n_211),
.C1(n_189),
.C2(n_207),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_196),
.C(n_182),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_305),
.B(n_217),
.CI(n_232),
.CON(n_307),
.SN(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_309),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_211),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.C(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_184),
.B1(n_207),
.B2(n_189),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_139),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_139),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.Y(n_320)
);


endmodule