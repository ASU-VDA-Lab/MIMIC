module fake_netlist_1_11381_n_655 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_655);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_655;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_599;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_48), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_56), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_3), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_50), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_62), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_66), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_64), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_77), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_30), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_76), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_69), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_54), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_45), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_5), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_14), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_60), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_35), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_47), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_57), .Y(n_112) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_25), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_27), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_5), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_114), .B(n_0), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_96), .B(n_0), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_81), .B(n_1), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_81), .B(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_79), .B(n_36), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_108), .A2(n_2), .B1(n_4), .B2(n_6), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_119), .B(n_2), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_119), .Y(n_132) );
BUFx8_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_108), .B(n_4), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_105), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_89), .B(n_7), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g145 ( .A1(n_116), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g147 ( .A1(n_89), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
AOI22x1_ASAP7_75t_SL g150 ( .A1(n_99), .A2(n_13), .B1(n_16), .B2(n_17), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_94), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_152) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_92), .A2(n_49), .B(n_20), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_78), .B(n_19), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_79), .B(n_19), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_142), .B(n_90), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_142), .B(n_90), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_124), .B(n_102), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_128), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_133), .B(n_103), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_121), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_123), .B(n_118), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_133), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_123), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_133), .B(n_84), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_122), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_135), .B(n_103), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_124), .B(n_117), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_155), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_126), .B(n_131), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_155), .B(n_93), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_126), .B(n_115), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_131), .B(n_100), .Y(n_184) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_127), .B(n_93), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_151), .B(n_80), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_150), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
BUFx6f_ASAP7_75t_SL g189 ( .A(n_127), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
INVx5_ASAP7_75t_L g191 ( .A(n_127), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_151), .B(n_149), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_120), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_132), .B(n_97), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_130), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_190), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_181), .B(n_130), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_166), .A2(n_150), .B1(n_145), .B2(n_147), .Y(n_201) );
INVxp67_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_198), .A2(n_125), .B1(n_143), .B2(n_129), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_198), .B(n_125), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_179), .A2(n_125), .B1(n_143), .B2(n_127), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_181), .B(n_143), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_179), .B(n_148), .Y(n_207) );
OAI22x1_ASAP7_75t_SL g208 ( .A1(n_187), .A2(n_140), .B1(n_129), .B2(n_152), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_175), .B(n_178), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_185), .A2(n_153), .B(n_149), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_196), .A2(n_104), .B(n_106), .C(n_132), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_159), .B(n_154), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_191), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_178), .B(n_88), .Y(n_216) );
O2A1O1Ixp5_ASAP7_75t_L g217 ( .A1(n_171), .A2(n_107), .B(n_112), .C(n_95), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_168), .A2(n_127), .B1(n_132), .B2(n_152), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
AND2x6_ASAP7_75t_SL g220 ( .A(n_160), .B(n_140), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_168), .B(n_88), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_168), .A2(n_92), .B1(n_113), .B2(n_111), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_168), .A2(n_113), .B1(n_109), .B2(n_98), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_176), .B(n_101), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_164), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_172), .A2(n_101), .B1(n_153), .B2(n_141), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_171), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_172), .B(n_173), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_172), .B(n_153), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_164), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_170), .B(n_153), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_172), .B(n_144), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g236 ( .A1(n_173), .A2(n_144), .B1(n_141), .B2(n_137), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_173), .B(n_144), .Y(n_237) );
AND2x6_ASAP7_75t_SL g238 ( .A(n_197), .B(n_144), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_183), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_173), .B(n_144), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_161), .B(n_141), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_171), .B(n_141), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_161), .B(n_141), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_182), .B(n_137), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_182), .B(n_137), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_186), .B(n_137), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_232), .A2(n_191), .B(n_180), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_199), .Y(n_252) );
INVx3_ASAP7_75t_SL g253 ( .A(n_230), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_209), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_200), .B(n_165), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_204), .B(n_174), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_204), .B(n_186), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_202), .B(n_191), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_231), .A2(n_191), .B(n_195), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_212), .A2(n_194), .B(n_193), .C(n_177), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_213), .B(n_184), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_216), .B(n_191), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_210), .A2(n_244), .B(n_205), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_230), .Y(n_264) );
NOR2x1_ASAP7_75t_R g265 ( .A(n_208), .B(n_191), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_219), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_206), .A2(n_194), .B(n_193), .C(n_169), .Y(n_268) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_243), .B(n_189), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_230), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_207), .A2(n_188), .B(n_169), .C(n_167), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g273 ( .A(n_201), .B(n_188), .C(n_169), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_215), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_224), .B(n_137), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_189), .B(n_188), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_SL g277 ( .A1(n_234), .A2(n_189), .B(n_167), .C(n_163), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_219), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_234), .B(n_21), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_218), .B(n_134), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_229), .A2(n_167), .B(n_163), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
CKINVDCx14_ASAP7_75t_R g285 ( .A(n_203), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_199), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_227), .A2(n_163), .B(n_162), .C(n_156), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_237), .A2(n_189), .B(n_162), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_203), .B(n_22), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_223), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_223), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_224), .B(n_134), .Y(n_292) );
O2A1O1Ixp5_ASAP7_75t_L g293 ( .A1(n_217), .A2(n_162), .B(n_156), .C(n_29), .Y(n_293) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_220), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_233), .A2(n_134), .B1(n_156), .B2(n_33), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_215), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_225), .B(n_134), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_SL g298 ( .A1(n_282), .A2(n_266), .B(n_278), .C(n_281), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_263), .A2(n_229), .B(n_246), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_294), .Y(n_300) );
NAND3x1_ASAP7_75t_L g301 ( .A(n_265), .B(n_208), .C(n_226), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_285), .A2(n_246), .B1(n_233), .B2(n_240), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_283), .A2(n_240), .B(n_239), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_254), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_251), .A2(n_241), .B(n_230), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_277), .A2(n_230), .B(n_214), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_276), .A2(n_214), .B(n_243), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_261), .A2(n_221), .B(n_239), .C(n_248), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_254), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
CKINVDCx6p67_ASAP7_75t_R g311 ( .A(n_294), .Y(n_311) );
AO21x1_ASAP7_75t_L g312 ( .A1(n_282), .A2(n_250), .B(n_249), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_266), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_247), .B(n_245), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_278), .B(n_248), .Y(n_315) );
AO31x2_ASAP7_75t_L g316 ( .A1(n_281), .A2(n_242), .A3(n_221), .B(n_236), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_288), .A2(n_228), .B(n_24), .Y(n_317) );
NOR4xp25_ASAP7_75t_L g318 ( .A(n_273), .B(n_23), .C(n_37), .D(n_39), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_SL g319 ( .A1(n_275), .A2(n_40), .B(n_42), .C(n_44), .Y(n_319) );
AO31x2_ASAP7_75t_L g320 ( .A1(n_292), .A2(n_228), .A3(n_51), .B(n_52), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_289), .A2(n_228), .B1(n_53), .B2(n_55), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_259), .A2(n_228), .B(n_58), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_284), .B(n_228), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_256), .B(n_46), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_296), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_297), .A2(n_61), .B(n_63), .C(n_65), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_257), .B(n_67), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_267), .A2(n_70), .B(n_71), .C(n_73), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_293), .A2(n_74), .B(n_75), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_267), .B(n_274), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_330), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_330), .Y(n_332) );
OAI21x1_ASAP7_75t_SL g333 ( .A1(n_303), .A2(n_274), .B(n_272), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_310), .A2(n_260), .B1(n_268), .B2(n_279), .C(n_272), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_302), .A2(n_279), .B1(n_258), .B2(n_262), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_298), .A2(n_280), .B(n_271), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_304), .A2(n_258), .B1(n_269), .B2(n_252), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_325), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_299), .A2(n_280), .B(n_295), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_313), .B(n_291), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
AOI211x1_ASAP7_75t_L g342 ( .A1(n_303), .A2(n_265), .B(n_258), .C(n_287), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_309), .B(n_253), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_314), .A2(n_264), .B(n_270), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_301), .B(n_258), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_327), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_299), .A2(n_270), .B1(n_264), .B2(n_290), .C(n_286), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_312), .A2(n_264), .B(n_270), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_329), .A2(n_253), .B(n_290), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_323), .B(n_253), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_317), .A2(n_252), .B(n_291), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_300), .A2(n_269), .B1(n_318), .B2(n_321), .C(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_311), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_336), .A2(n_326), .B(n_319), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_345), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_341), .B(n_323), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_342), .B(n_321), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_333), .A2(n_306), .B(n_305), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_331), .B(n_320), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_341), .B(n_316), .Y(n_364) );
OA21x2_ASAP7_75t_L g365 ( .A1(n_346), .A2(n_322), .B(n_307), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_346), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_354), .A2(n_320), .B(n_316), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_331), .B(n_320), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_343), .B(n_316), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_332), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_338), .A2(n_269), .B1(n_328), .B2(n_334), .C(n_355), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_333), .A2(n_350), .B(n_352), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_353), .Y(n_375) );
AO21x1_ASAP7_75t_SL g376 ( .A1(n_343), .A2(n_356), .B(n_351), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_344), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_347), .B(n_351), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_354), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_356), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_357), .Y(n_383) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_339), .B(n_340), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_352), .A2(n_339), .B(n_349), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_363), .B(n_339), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_367), .A2(n_339), .B(n_337), .Y(n_389) );
OA21x2_ASAP7_75t_L g390 ( .A1(n_367), .A2(n_335), .B(n_381), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_382), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_382), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_364), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_364), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_378), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_363), .B(n_368), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_361), .A2(n_359), .B1(n_373), .B2(n_375), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
BUFx5_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_368), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_380), .B(n_372), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_368), .B(n_379), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_361), .A2(n_375), .B1(n_386), .B2(n_385), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
OR2x6_ASAP7_75t_L g413 ( .A(n_361), .B(n_380), .Y(n_413) );
AO21x2_ASAP7_75t_L g414 ( .A1(n_381), .A2(n_387), .B(n_358), .Y(n_414) );
INVx5_ASAP7_75t_SL g415 ( .A(n_361), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_377), .B(n_379), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_377), .B(n_360), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_360), .B(n_369), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
INVx4_ASAP7_75t_L g420 ( .A(n_361), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_374), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_366), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_374), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_374), .B(n_387), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_362), .B(n_366), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_387), .B(n_376), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_362), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_366), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_362), .B(n_381), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_399), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_410), .B(n_376), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_418), .B(n_383), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_400), .A2(n_385), .B(n_386), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_430), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_398), .B(n_358), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_418), .B(n_365), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_410), .B(n_365), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_395), .B(n_365), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_399), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_410), .B(n_365), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_408), .B(n_358), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_398), .B(n_426), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_403), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_393), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_393), .B(n_394), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_393), .B(n_397), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_408), .B(n_417), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_404), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_417), .B(n_392), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_417), .B(n_392), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_406), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_394), .B(n_396), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
BUFx2_ASAP7_75t_SL g459 ( .A(n_406), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_394), .B(n_396), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_391), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_396), .B(n_397), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_397), .B(n_421), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_421), .B(n_424), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_400), .B(n_401), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_426), .B(n_407), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_416), .B(n_402), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_401), .B(n_405), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_421), .B(n_424), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_420), .B(n_419), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_416), .B(n_424), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_426), .B(n_407), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_405), .B(n_413), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_425), .B(n_416), .Y(n_475) );
NAND3xp33_ASAP7_75t_SL g476 ( .A(n_411), .B(n_428), .C(n_420), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
NAND2xp33_ASAP7_75t_L g479 ( .A(n_406), .B(n_427), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_425), .B(n_388), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_425), .B(n_419), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_388), .B(n_413), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_388), .B(n_413), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_406), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_413), .B(n_420), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_427), .B(n_415), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_467), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_480), .B(n_465), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_472), .B(n_413), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_475), .B(n_427), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_441), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_452), .Y(n_495) );
NAND2xp33_ASAP7_75t_L g496 ( .A(n_456), .B(n_406), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_433), .B(n_420), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_475), .B(n_415), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_456), .Y(n_500) );
NAND3x1_ASAP7_75t_L g501 ( .A(n_432), .B(n_415), .C(n_413), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_467), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_451), .B(n_415), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_468), .B(n_426), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_441), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_445), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_480), .B(n_406), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_465), .B(n_406), .Y(n_508) );
XNOR2xp5_ASAP7_75t_L g509 ( .A(n_432), .B(n_426), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_454), .B(n_415), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_470), .B(n_415), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_435), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_471), .B(n_423), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_470), .B(n_406), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_482), .B(n_406), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_447), .B(n_406), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_455), .B(n_406), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_447), .B(n_390), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_469), .B(n_390), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_466), .B(n_390), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_459), .A2(n_423), .B1(n_390), .B2(n_389), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_483), .B(n_390), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_464), .B(n_389), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_464), .B(n_389), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_440), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_466), .B(n_423), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_444), .B(n_389), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_469), .B(n_429), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_444), .B(n_414), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_445), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_444), .B(n_414), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_485), .B(n_409), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
OAI332xp33_ASAP7_75t_L g535 ( .A1(n_443), .A2(n_409), .A3(n_412), .B1(n_414), .B2(n_422), .B3(n_429), .C1(n_438), .C2(n_478), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_448), .B(n_429), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_449), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_453), .B(n_414), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_483), .B(n_409), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_453), .B(n_412), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_458), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_439), .B(n_412), .Y(n_543) );
NOR2x1p5_ASAP7_75t_L g544 ( .A(n_476), .B(n_474), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_490), .B(n_484), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_498), .A2(n_484), .B1(n_439), .B2(n_442), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_490), .B(n_538), .Y(n_547) );
NAND2xp33_ASAP7_75t_SL g548 ( .A(n_544), .B(n_474), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_500), .B(n_471), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_512), .A2(n_434), .B(n_479), .C(n_485), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_488), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_442), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_504), .B(n_458), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_513), .B(n_467), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_500), .B(n_434), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_518), .B(n_462), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_491), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_535), .B(n_462), .C(n_440), .Y(n_558) );
OAI22xp33_ASAP7_75t_SL g559 ( .A1(n_489), .A2(n_487), .B1(n_473), .B2(n_467), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_518), .B(n_457), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_494), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_507), .Y(n_564) );
AOI32xp33_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_473), .A3(n_486), .B1(n_437), .B2(n_481), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_506), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_531), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_493), .B(n_457), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_509), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_537), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_508), .B(n_459), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_522), .Y(n_574) );
NOR3xp33_ASAP7_75t_L g575 ( .A(n_520), .B(n_481), .C(n_436), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_486), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_543), .B(n_450), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_489), .B(n_473), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_450), .Y(n_581) );
XOR2xp5_ASAP7_75t_L g582 ( .A(n_503), .B(n_437), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_495), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_517), .B(n_536), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_542), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_542), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_567), .B(n_523), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_558), .B(n_539), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_556), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_567), .B(n_519), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_548), .A2(n_498), .B1(n_525), .B2(n_524), .C1(n_496), .C2(n_528), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_577), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_577), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_549), .B(n_513), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_557), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_562), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_558), .B(n_543), .Y(n_599) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_555), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_547), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_563), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_555), .A2(n_533), .B(n_513), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_566), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_575), .B(n_530), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_571), .A2(n_548), .B1(n_575), .B2(n_546), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g607 ( .A1(n_559), .A2(n_527), .B(n_532), .C(n_530), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_565), .B(n_489), .Y(n_609) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_583), .Y(n_610) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_549), .A2(n_502), .B(n_514), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_569), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_560), .B(n_529), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_606), .A2(n_550), .B1(n_554), .B2(n_553), .C(n_582), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_609), .B(n_564), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_589), .A2(n_561), .B1(n_552), .B2(n_572), .C(n_545), .Y(n_616) );
XNOR2x1_ASAP7_75t_L g617 ( .A(n_599), .B(n_554), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_607), .A2(n_501), .B1(n_580), .B2(n_502), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_589), .B(n_584), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g620 ( .A1(n_611), .A2(n_502), .B(n_573), .C(n_521), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_594), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_600), .A2(n_578), .A3(n_579), .B1(n_580), .B2(n_514), .C1(n_528), .C2(n_532), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_605), .A2(n_580), .B1(n_527), .B2(n_585), .C(n_586), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_591), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_592), .A2(n_533), .B(n_587), .Y(n_625) );
AOI21xp5_ASAP7_75t_SL g626 ( .A1(n_603), .A2(n_501), .B(n_511), .Y(n_626) );
OAI32xp33_ASAP7_75t_L g627 ( .A1(n_596), .A2(n_570), .A3(n_581), .B1(n_492), .B2(n_499), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_595), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_593), .A2(n_583), .B1(n_574), .B2(n_576), .C1(n_437), .C2(n_516), .Y(n_629) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_614), .A2(n_592), .B(n_612), .Y(n_630) );
NOR2xp33_ASAP7_75t_R g631 ( .A(n_624), .B(n_601), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_618), .A2(n_590), .B1(n_604), .B2(n_608), .C(n_602), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_619), .A2(n_596), .B1(n_588), .B2(n_598), .Y(n_633) );
AOI211xp5_ASAP7_75t_SL g634 ( .A1(n_626), .A2(n_610), .B(n_510), .C(n_597), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_615), .A2(n_437), .B1(n_473), .B2(n_516), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_620), .A2(n_613), .B(n_540), .C(n_576), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_616), .B(n_574), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_625), .A2(n_541), .B(n_497), .C(n_446), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g639 ( .A(n_634), .B(n_629), .C(n_622), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_632), .B(n_627), .C(n_623), .Y(n_640) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_630), .A2(n_629), .B(n_621), .C(n_628), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_637), .B(n_617), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_638), .B(n_497), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_641), .A2(n_636), .B(n_633), .Y(n_644) );
OR5x1_ASAP7_75t_L g645 ( .A(n_639), .B(n_631), .C(n_635), .D(n_446), .E(n_436), .Y(n_645) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_642), .B(n_448), .C(n_463), .D(n_461), .E(n_460), .Y(n_646) );
AND2x2_ASAP7_75t_SL g647 ( .A(n_645), .B(n_640), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_644), .Y(n_648) );
OAI22xp5_ASAP7_75t_SL g649 ( .A1(n_648), .A2(n_643), .B1(n_646), .B2(n_446), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_648), .Y(n_650) );
AOI22x1_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_647), .B1(n_436), .B2(n_460), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
OAI21x1_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_647), .B(n_649), .Y(n_653) );
OAI32xp33_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_460), .A3(n_477), .B1(n_422), .B2(n_463), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_477), .B1(n_461), .B2(n_422), .Y(n_655) );
endmodule