module fake_jpeg_18092_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_11),
.B(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_23),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_4),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_81),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_64),
.B1(n_62),
.B2(n_51),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_51),
.B1(n_58),
.B2(n_73),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_85),
.B1(n_92),
.B2(n_88),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_61),
.C(n_68),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_72),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_71),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_54),
.B1(n_50),
.B2(n_59),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_94),
.B(n_102),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_88),
.B1(n_70),
.B2(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_52),
.B1(n_48),
.B2(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_52),
.B1(n_63),
.B2(n_55),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_111),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_69),
.B1(n_60),
.B2(n_48),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_20),
.B(n_21),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_112),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_57),
.B(n_56),
.C(n_74),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_118),
.B1(n_121),
.B2(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_47),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_8),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_130),
.B1(n_111),
.B2(n_34),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_17),
.C(n_19),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_133),
.C(n_108),
.Y(n_135)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_24),
.B(n_27),
.C(n_28),
.D(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_30),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_137),
.Y(n_144)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_129),
.B1(n_133),
.B2(n_36),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_131),
.B1(n_132),
.B2(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_139),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_140),
.Y(n_157)
);

OAI321xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_149),
.A3(n_143),
.B1(n_144),
.B2(n_141),
.C(n_135),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_143),
.C(n_35),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_41),
.Y(n_160)
);


endmodule