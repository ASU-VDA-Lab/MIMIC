module real_jpeg_528_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_45),
.B1(n_67),
.B2(n_69),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_41),
.B1(n_67),
.B2(n_69),
.Y(n_181)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_4),
.A2(n_67),
.B1(n_69),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_42),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_30),
.B(n_85),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_48),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_39),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_64),
.C(n_67),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_5),
.B(n_78),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_108),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_67),
.B1(n_69),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_6),
.Y(n_104)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_37),
.B1(n_39),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_57),
.B1(n_67),
.B2(n_69),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_67),
.B1(n_69),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_12),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_74),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_97),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_97),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_13),
.A2(n_67),
.B1(n_69),
.B2(n_97),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_14),
.A2(n_27),
.B1(n_67),
.B2(n_69),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_16),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_16),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_16),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_16),
.A2(n_37),
.B1(n_39),
.B2(n_71),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_131),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_110),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_22),
.B(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_99),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_23),
.B(n_99),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_58),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_25),
.B(n_43),
.C(n_58),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_42),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_28),
.A2(n_34),
.A3(n_39),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_33),
.B(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_36),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_36),
.A2(n_95),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_36),
.A2(n_95),
.B1(n_96),
.B2(n_165),
.Y(n_164)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_39),
.B1(n_52),
.B2(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_37),
.B(n_153),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_39),
.A2(n_50),
.A3(n_52),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_56),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_92),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_47),
.A2(n_92),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_47),
.A2(n_91),
.B1(n_92),
.B2(n_139),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_47),
.A2(n_92),
.B1(n_138),
.B2(n_186),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AO22x2_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_49),
.B(n_54),
.Y(n_154)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_50),
.B(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_56),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_72),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_59),
.B(n_72),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_66),
.B2(n_70),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_61),
.A2(n_66),
.B1(n_148),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_62),
.A2(n_107),
.B1(n_108),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_62),
.A2(n_108),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_62),
.A2(n_108),
.B1(n_149),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_62),
.A2(n_108),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_62),
.A2(n_108),
.B1(n_177),
.B2(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_67),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_80),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_77),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_75),
.A2(n_77),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_75),
.A2(n_77),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_78),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_78),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_76),
.A2(n_78),
.B1(n_88),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_76),
.A2(n_78),
.B1(n_157),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_76),
.A2(n_78),
.B1(n_153),
.B2(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_76),
.A2(n_78),
.B1(n_207),
.B2(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_82),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.C(n_94),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_83),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_87),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_90),
.B(n_94),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_109),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_129),
.B2(n_130),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

AOI31xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_227),
.A3(n_236),
.B(n_240),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_172),
.B(n_226),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_159),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_159),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.C(n_150),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_136),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_141),
.C(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_146),
.B(n_150),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_167),
.C(n_171),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_221),
.B(n_225),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_190),
.B(n_220),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_182),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_179),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_185),
.C(n_188),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_201),
.B(n_219),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_213),
.B(n_218),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_212),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_224),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_235),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);


endmodule