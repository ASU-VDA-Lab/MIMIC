module fake_jpeg_28472_n_453 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_83),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_38),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_43),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_98),
.Y(n_155)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_48),
.B1(n_46),
.B2(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_41),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_49),
.C(n_28),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_103),
.B(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_31),
.B1(n_23),
.B2(n_45),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_3),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_3),
.B(n_4),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_49),
.B1(n_45),
.B2(n_44),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_151),
.B1(n_154),
.B2(n_47),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_71),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_84),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_58),
.A2(n_48),
.B1(n_46),
.B2(n_34),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_152),
.B1(n_50),
.B2(n_73),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_24),
.B1(n_47),
.B2(n_25),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_83),
.A2(n_48),
.B1(n_46),
.B2(n_34),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_63),
.A2(n_23),
.B1(n_44),
.B2(n_43),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_123),
.B(n_152),
.Y(n_217)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_101),
.A2(n_85),
.B1(n_48),
.B2(n_34),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_36),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_169),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_36),
.B(n_40),
.C(n_28),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_166),
.B(n_188),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_40),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_25),
.B(n_24),
.C(n_46),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_181),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_130),
.Y(n_173)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_66),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_187),
.Y(n_211)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_177),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_67),
.B1(n_76),
.B2(n_70),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_186),
.B1(n_197),
.B2(n_199),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_96),
.B1(n_93),
.B2(n_91),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_113),
.A2(n_87),
.B1(n_80),
.B2(n_78),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_77),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_190),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_150),
.B(n_4),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_7),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_138),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_8),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_191),
.B1(n_183),
.B2(n_170),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_161),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_169),
.C(n_165),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_191),
.C(n_160),
.Y(n_253)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_183),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_253),
.C(n_248),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_171),
.B1(n_157),
.B2(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_256),
.Y(n_279)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_205),
.B(n_166),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_248),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_257),
.B1(n_262),
.B2(n_210),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_198),
.C(n_196),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_252),
.B(n_265),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_253),
.B(n_179),
.Y(n_290)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_214),
.A2(n_181),
.B(n_187),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_255),
.A2(n_266),
.B(n_174),
.Y(n_294)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_211),
.A2(n_128),
.B1(n_197),
.B2(n_126),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_211),
.A2(n_236),
.B1(n_208),
.B2(n_226),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_270),
.B1(n_277),
.B2(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_217),
.B1(n_223),
.B2(n_229),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_227),
.C(n_205),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_274),
.C(n_293),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_210),
.B(n_216),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_275),
.B(n_281),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_229),
.B(n_206),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_216),
.B1(n_115),
.B2(n_159),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_215),
.B(n_202),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_228),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_289),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_215),
.B(n_207),
.C(n_234),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_283),
.B(n_294),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_207),
.B1(n_200),
.B2(n_143),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_168),
.B1(n_132),
.B2(n_107),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_291),
.B1(n_285),
.B2(n_209),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_163),
.B(n_233),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_193),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_242),
.A2(n_132),
.B1(n_143),
.B2(n_107),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_233),
.C(n_213),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_242),
.B1(n_238),
.B2(n_224),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_315),
.B1(n_320),
.B2(n_267),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

AO22x1_ASAP7_75t_SL g297 ( 
.A1(n_279),
.A2(n_206),
.B1(n_241),
.B2(n_212),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_213),
.Y(n_301)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_303),
.B(n_158),
.Y(n_337)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_224),
.B1(n_209),
.B2(n_222),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_305),
.A2(n_306),
.B1(n_291),
.B2(n_292),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_276),
.A2(n_264),
.B1(n_206),
.B2(n_220),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_311),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_194),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_276),
.B(n_277),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_316),
.B(n_178),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_282),
.B1(n_269),
.B2(n_294),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_317),
.A2(n_318),
.B1(n_284),
.B2(n_271),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_222),
.B1(n_104),
.B2(n_149),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_225),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_319),
.Y(n_326)
);

OAI22x1_ASAP7_75t_L g320 ( 
.A1(n_280),
.A2(n_273),
.B1(n_286),
.B2(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_289),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_332),
.B1(n_342),
.B2(n_190),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_274),
.C(n_290),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_343),
.C(n_298),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_290),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_333),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_286),
.B(n_293),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_192),
.B(n_173),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_219),
.B(n_292),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_305),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_335),
.A2(n_339),
.B1(n_315),
.B2(n_318),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_288),
.B1(n_149),
.B2(n_146),
.Y(n_336)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_299),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_301),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_338),
.B(n_341),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_288),
.B1(n_219),
.B2(n_188),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_307),
.A2(n_250),
.B1(n_230),
.B2(n_182),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_225),
.C(n_175),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_136),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_297),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_298),
.CI(n_309),
.CON(n_350),
.SN(n_350)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_351),
.B(n_363),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_353),
.A2(n_361),
.B1(n_342),
.B2(n_348),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_356),
.C(n_364),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_309),
.C(n_319),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_297),
.Y(n_358)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_310),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_369),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_250),
.B1(n_173),
.B2(n_167),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_330),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_334),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_195),
.C(n_189),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_365),
.A2(n_335),
.B1(n_340),
.B2(n_344),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_201),
.C(n_134),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_332),
.C(n_333),
.Y(n_375)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_239),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_328),
.B1(n_347),
.B2(n_339),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_373),
.A2(n_353),
.B1(n_362),
.B2(n_370),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_379),
.C(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_331),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_350),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_346),
.C(n_330),
.Y(n_379)
);

AOI31xp33_ASAP7_75t_L g380 ( 
.A1(n_370),
.A2(n_348),
.A3(n_323),
.B(n_325),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_380),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_384),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_382),
.A2(n_344),
.B1(n_368),
.B2(n_369),
.Y(n_404)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_352),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_364),
.C(n_359),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_367),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_391),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_387),
.B(n_374),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_397),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_375),
.C(n_385),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_401),
.C(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_366),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_389),
.A2(n_349),
.B(n_358),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_404),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_365),
.C(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_402),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_350),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_386),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_377),
.B(n_347),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_405),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_392),
.A2(n_400),
.B(n_403),
.Y(n_406)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_406),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_372),
.C(n_384),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_382),
.C(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_410),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_114),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_328),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_418),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_373),
.C(n_389),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_139),
.C(n_137),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_361),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_398),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_421),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_396),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_396),
.B(n_180),
.Y(n_424)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_425),
.B(n_426),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_148),
.B1(n_118),
.B2(n_122),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_416),
.A2(n_114),
.B1(n_118),
.B2(n_11),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_427),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_429),
.A2(n_431),
.B(n_414),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g439 ( 
.A(n_430),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_412),
.B(n_9),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_434),
.B(n_425),
.Y(n_440)
);

AOI21xp33_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_428),
.B(n_423),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_435),
.A2(n_438),
.B(n_430),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_423),
.A2(n_417),
.B(n_418),
.Y(n_438)
);

A2O1A1O1Ixp25_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_436),
.B(n_439),
.C(n_12),
.D(n_13),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_417),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_SL g447 ( 
.A1(n_441),
.A2(n_442),
.B(n_444),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_437),
.Y(n_443)
);

OAI21x1_ASAP7_75t_SL g446 ( 
.A1(n_443),
.A2(n_10),
.B(n_11),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_426),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_446),
.B(n_13),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_449),
.A2(n_447),
.B(n_14),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_448),
.B(n_14),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_14),
.Y(n_453)
);


endmodule