module fake_jpeg_19318_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

AND2x6_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_19),
.B(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_20),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_6),
.B1(n_2),
.B2(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_2),
.B1(n_6),
.B2(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_28),
.C(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_28),
.B1(n_16),
.B2(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_14),
.B1(n_29),
.B2(n_35),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_34),
.Y(n_39)
);

AOI21x1_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_41),
.B(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_40)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_24),
.C(n_25),
.Y(n_41)
);

OAI21x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_37),
.B(n_14),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_39),
.B(n_14),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.C(n_45),
.Y(n_47)
);


endmodule