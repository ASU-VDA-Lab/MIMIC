module fake_jpeg_5162_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_9),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_34),
.B(n_28),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_56),
.Y(n_90)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_18),
.B1(n_46),
.B2(n_42),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_78),
.B1(n_65),
.B2(n_71),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_45),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_42),
.B1(n_23),
.B2(n_45),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_32),
.B1(n_31),
.B2(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_43),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_43),
.B1(n_46),
.B2(n_32),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_35),
.C(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_62),
.B1(n_68),
.B2(n_59),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_84),
.B(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_113),
.Y(n_147)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_118),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_34),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_120),
.Y(n_153)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_67),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_58),
.B1(n_57),
.B2(n_70),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_125),
.C(n_128),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_53),
.C(n_51),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_69),
.CI(n_50),
.CON(n_127),
.SN(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_131),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_56),
.C(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_129),
.Y(n_135)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_33),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_100),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_157),
.B(n_30),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_126),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_86),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_82),
.B1(n_83),
.B2(n_21),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_84),
.Y(n_145)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_127),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_34),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_165),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_115),
.B1(n_127),
.B2(n_117),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_164),
.B1(n_184),
.B2(n_154),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_115),
.A3(n_104),
.B1(n_114),
.B2(n_112),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_184),
.Y(n_210)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_128),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_170),
.B(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_82),
.B1(n_83),
.B2(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_35),
.B(n_21),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_146),
.B1(n_141),
.B2(n_136),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_116),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_123),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_141),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_34),
.B(n_28),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_148),
.B1(n_140),
.B2(n_133),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_193),
.B1(n_144),
.B2(n_152),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_149),
.C(n_138),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_198),
.C(n_212),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_163),
.B1(n_157),
.B2(n_166),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_149),
.C(n_138),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_170),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_157),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_144),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_159),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_150),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_136),
.C(n_146),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_214),
.C(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_165),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_220),
.B(n_224),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_169),
.B1(n_158),
.B2(n_126),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_231),
.B1(n_233),
.B2(n_17),
.Y(n_258)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_202),
.B1(n_207),
.B2(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_235),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_148),
.B1(n_140),
.B2(n_113),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_28),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_156),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_209),
.B(n_190),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_215),
.A2(n_192),
.B(n_193),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_257),
.B1(n_213),
.B2(n_221),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_198),
.B1(n_192),
.B2(n_197),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_28),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_209),
.B1(n_188),
.B2(n_150),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_229),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_135),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_135),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_99),
.B(n_30),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_0),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_237),
.C(n_219),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_267),
.C(n_272),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_260),
.B(n_253),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_243),
.B1(n_239),
.B2(n_240),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_156),
.C(n_120),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_110),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_279),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_280),
.B1(n_250),
.B2(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_72),
.C(n_26),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_26),
.C(n_25),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.C(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_30),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_29),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_265),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_240),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_287),
.B(n_290),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_283),
.A2(n_289),
.B1(n_296),
.B2(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_260),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_294),
.B(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_247),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_291),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_245),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_25),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_241),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_253),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_262),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_266),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_290),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_267),
.C(n_257),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_309),
.C(n_1),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_278),
.B1(n_255),
.B2(n_242),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_241),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_29),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_289),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_315),
.B(n_319),
.Y(n_327)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_17),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_320),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_0),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_0),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_1),
.C(n_5),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_299),
.B1(n_309),
.B2(n_298),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_325),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_307),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_314),
.A3(n_316),
.B1(n_321),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_324),
.A2(n_326),
.B(n_6),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_318),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_311),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_7),
.B(n_8),
.C(n_10),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_333),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_334),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_11),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_329),
.A3(n_331),
.B1(n_328),
.B2(n_324),
.C1(n_16),
.C2(n_14),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_336),
.B(n_12),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_12),
.C(n_14),
.Y(n_340)
);

NAND4xp25_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_12),
.C(n_14),
.D(n_16),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_16),
.Y(n_342)
);


endmodule