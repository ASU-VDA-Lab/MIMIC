module fake_netlist_6_2584_n_1882 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1882);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1882;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g197 ( 
.A(n_42),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_69),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_63),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_78),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_106),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_1),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_88),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_64),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_14),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_85),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_114),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_134),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_83),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_111),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_23),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_119),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_72),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_2),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_39),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_133),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_172),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_97),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_93),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_149),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_109),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_34),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_26),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_18),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_22),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_59),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_62),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_91),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_31),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_195),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_26),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_73),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_171),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_13),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_96),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_38),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_107),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_84),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_44),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_117),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_58),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_176),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_53),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_65),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_81),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_103),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_108),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_92),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_140),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_55),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_174),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_170),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_173),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_180),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_57),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_82),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_175),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_30),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_113),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_13),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_21),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_39),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_28),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_87),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_50),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_148),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_152),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_56),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_20),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_161),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_100),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_51),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_24),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_32),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_25),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_123),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_144),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_168),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_68),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_55),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_48),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_50),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_44),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_188),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_128),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_186),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_179),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_190),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_167),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_71),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_112),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_76),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_157),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_131),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_135),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_46),
.Y(n_345)
);

BUFx2_ASAP7_75t_R g346 ( 
.A(n_5),
.Y(n_346)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_80),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_193),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_30),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_159),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_23),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_125),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_162),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_14),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_102),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_15),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_153),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_67),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_124),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_156),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_52),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_141),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_56),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_118),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_138),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_145),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_54),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_25),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_126),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_74),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_181),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_8),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_61),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_60),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_165),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_89),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_19),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_27),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_60),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_51),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_189),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_43),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_191),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_35),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_187),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_0),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_130),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_9),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_31),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_121),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_197),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_202),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_200),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_257),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_202),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_207),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_368),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_207),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_209),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_209),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_214),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_201),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_210),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_199),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_206),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_240),
.B(n_3),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_216),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_232),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_212),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_257),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_245),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_268),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_258),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_296),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_208),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_217),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_301),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_366),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_219),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_208),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_224),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_218),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_214),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_219),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_225),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_239),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_239),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_233),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_280),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_247),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_236),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_198),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_203),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_237),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_247),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_254),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_255),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_241),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_255),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_270),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_218),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_199),
.B(n_3),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_204),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_223),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_205),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_221),
.B(n_4),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_250),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_270),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_211),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_213),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_275),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_275),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_252),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_251),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_256),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_261),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_252),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_220),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_222),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_262),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_277),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_277),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_283),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_267),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_328),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_283),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_291),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_291),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_221),
.B(n_4),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_293),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_274),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_279),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_282),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_328),
.B(n_334),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_285),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_226),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_293),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_288),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_R g484 ( 
.A(n_228),
.B(n_192),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_292),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_334),
.B(n_6),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_230),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_231),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_297),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_234),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_297),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_298),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_215),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_406),
.B(n_344),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_435),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_436),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_448),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_394),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_447),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_449),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_453),
.Y(n_512)
);

BUFx8_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_454),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_344),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_397),
.B(n_229),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_399),
.B(n_361),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_458),
.B(n_361),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_400),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_463),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_404),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_464),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_229),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_415),
.B(n_260),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_481),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_488),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_432),
.B(n_235),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_398),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_260),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_462),
.B(n_266),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_438),
.A2(n_327),
.B(n_284),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_440),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_350),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_452),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_266),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_490),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_SL g548 ( 
.A(n_426),
.B(n_271),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_405),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_470),
.B(n_353),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_409),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_457),
.B(n_353),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_409),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_456),
.B(n_358),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_465),
.B(n_350),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_466),
.A2(n_327),
.B(n_284),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_468),
.B(n_358),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g561 ( 
.A(n_417),
.B(n_333),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_418),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_418),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_407),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_428),
.B(n_238),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_509),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_515),
.A2(n_486),
.B1(n_446),
.B2(n_243),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_509),
.Y(n_576)
);

BUFx4f_ASAP7_75t_L g577 ( 
.A(n_546),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_573),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_503),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_554),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_569),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_497),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_510),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_557),
.B(n_431),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_515),
.B(n_402),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_569),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_497),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_494),
.A2(n_243),
.B1(n_265),
.B2(n_215),
.Y(n_590)
);

AND2x2_ASAP7_75t_SL g591 ( 
.A(n_494),
.B(n_333),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_546),
.B(n_431),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_518),
.A2(n_307),
.B1(n_345),
.B2(n_265),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_518),
.A2(n_345),
.B1(n_354),
.B2(n_307),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_546),
.B(n_434),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_538),
.B(n_469),
.C(n_437),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_511),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_525),
.B(n_434),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_500),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_550),
.B(n_465),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_548),
.A2(n_477),
.B1(n_451),
.B2(n_459),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_513),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_560),
.B(n_338),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_506),
.Y(n_606)
);

BUFx4f_ASAP7_75t_L g607 ( 
.A(n_560),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_516),
.B(n_338),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_569),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_513),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_528),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_517),
.B(n_487),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_517),
.A2(n_354),
.B1(n_385),
.B2(n_324),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_534),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_526),
.B(n_477),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_530),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_540),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_516),
.B(n_223),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_513),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_551),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_551),
.B(n_442),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_516),
.B(n_298),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_516),
.B(n_223),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_524),
.B(n_304),
.Y(n_634)
);

INVx4_ASAP7_75t_SL g635 ( 
.A(n_569),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_524),
.A2(n_385),
.B1(n_271),
.B2(n_324),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_535),
.B(n_451),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_507),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_498),
.B(n_395),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_541),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_564),
.B(n_459),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_552),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_524),
.B(n_223),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_570),
.B(n_460),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_524),
.B(n_223),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_564),
.B(n_460),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_564),
.B(n_461),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_571),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_537),
.B(n_382),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_537),
.B(n_304),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_555),
.B(n_346),
.Y(n_654)
);

OAI21xp33_ASAP7_75t_SL g655 ( 
.A1(n_539),
.A2(n_474),
.B(n_450),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_507),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_498),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_537),
.B(n_318),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_542),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_519),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_537),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_535),
.B(n_461),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_535),
.B(n_476),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_571),
.B(n_476),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_478),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_562),
.B(n_478),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_565),
.B(n_480),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_480),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_545),
.B(n_318),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_513),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_495),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_545),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_553),
.Y(n_674)
);

INVx4_ASAP7_75t_SL g675 ( 
.A(n_571),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_499),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_506),
.B(n_483),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_519),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_519),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_553),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_522),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_559),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_559),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_558),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_543),
.B(n_382),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_543),
.B(n_412),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_572),
.A2(n_381),
.B1(n_387),
.B2(n_312),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_563),
.B(n_483),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_485),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_566),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_520),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx4_ASAP7_75t_SL g694 ( 
.A(n_568),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_520),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_568),
.A2(n_281),
.B1(n_330),
.B2(n_269),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_572),
.B(n_242),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_520),
.B(n_244),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_531),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_504),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_531),
.B(n_382),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_533),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_558),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_533),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_533),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_536),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_536),
.B(n_382),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_536),
.A2(n_281),
.B1(n_330),
.B2(n_349),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_544),
.B(n_423),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_544),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_544),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_496),
.B(n_325),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_496),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_502),
.B(n_425),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_580),
.B(n_303),
.Y(n_715)
);

O2A1O1Ixp5_ASAP7_75t_L g716 ( 
.A1(n_620),
.A2(n_629),
.B(n_648),
.C(n_646),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_602),
.B(n_305),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_613),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_591),
.A2(n_410),
.B1(n_421),
.B2(n_420),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_602),
.B(n_309),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_577),
.B(n_382),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_585),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_657),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_666),
.B(n_325),
.Y(n_725)
);

AND3x1_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_246),
.C(n_227),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_313),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_591),
.A2(n_413),
.B1(n_419),
.B2(n_416),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_575),
.B(n_445),
.C(n_321),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_625),
.B(n_505),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_587),
.B(n_317),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_666),
.A2(n_414),
.B1(n_302),
.B2(n_388),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_607),
.A2(n_342),
.B1(n_341),
.B2(n_343),
.Y(n_734)
);

O2A1O1Ixp5_ASAP7_75t_L g735 ( 
.A1(n_620),
.A2(n_341),
.B(n_377),
.C(n_352),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_587),
.B(n_322),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_618),
.B(n_512),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_577),
.B(n_514),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_599),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_590),
.A2(n_294),
.B1(n_320),
.B2(n_316),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_661),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_590),
.A2(n_594),
.B1(n_593),
.B2(n_614),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_607),
.B(n_521),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_669),
.B(n_523),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_608),
.A2(n_263),
.B(n_349),
.C(n_248),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_695),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_695),
.B(n_658),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_713),
.B(n_665),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_592),
.B(n_527),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_612),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_615),
.B(n_372),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_616),
.B(n_372),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_700),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_619),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_689),
.B(n_690),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_595),
.B(n_529),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_632),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_641),
.B(n_642),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_679),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_660),
.B(n_376),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_617),
.A2(n_286),
.B1(n_249),
.B2(n_384),
.Y(n_764)
);

AND2x2_ASAP7_75t_SL g765 ( 
.A(n_593),
.B(n_376),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_643),
.B(n_547),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_673),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_674),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_617),
.A2(n_278),
.B1(n_253),
.B2(n_259),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_681),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_680),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_594),
.A2(n_227),
.B1(n_246),
.B2(n_248),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_683),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_649),
.B(n_484),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_693),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_650),
.B(n_272),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_687),
.B(n_640),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_684),
.B(n_377),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_650),
.B(n_273),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_638),
.B(n_386),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_663),
.B(n_664),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_709),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_299),
.B1(n_264),
.B2(n_269),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_634),
.B(n_508),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_705),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_676),
.B(n_685),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_508),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_689),
.B(n_331),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_690),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_682),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_634),
.B(n_287),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_688),
.A2(n_323),
.B1(n_308),
.B2(n_300),
.C(n_294),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_678),
.A2(n_264),
.B1(n_383),
.B2(n_375),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_574),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_578),
.B(n_289),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_634),
.B(n_290),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_653),
.B(n_380),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_667),
.B(n_230),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_598),
.B(n_332),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_574),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_624),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_702),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_L g805 ( 
.A1(n_696),
.A2(n_329),
.B1(n_360),
.B2(n_383),
.C(n_320),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_576),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_L g807 ( 
.A1(n_603),
.A2(n_360),
.B1(n_329),
.B2(n_364),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_704),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_697),
.B(n_351),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_668),
.B(n_624),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_703),
.A2(n_375),
.B1(n_276),
.B2(n_299),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_676),
.B(n_295),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_653),
.B(n_310),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_653),
.B(n_311),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_698),
.B(n_356),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_714),
.B(n_362),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_582),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_618),
.B(n_314),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_627),
.B(n_315),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_711),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_703),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_645),
.B(n_319),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_677),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_706),
.B(n_655),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_714),
.B(n_369),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_706),
.B(n_326),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_706),
.B(n_335),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_706),
.B(n_336),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_636),
.B(n_337),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_640),
.B(n_230),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_671),
.B(n_339),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_640),
.B(n_373),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_608),
.B(n_340),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_611),
.Y(n_834)
);

INVx8_ASAP7_75t_L g835 ( 
.A(n_677),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_626),
.B(n_230),
.Y(n_836)
);

AND2x2_ASAP7_75t_SL g837 ( 
.A(n_654),
.B(n_276),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_712),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_636),
.B(n_626),
.Y(n_839)
);

BUFx6f_ASAP7_75t_SL g840 ( 
.A(n_700),
.Y(n_840)
);

BUFx5_ASAP7_75t_L g841 ( 
.A(n_627),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_606),
.B(n_348),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_712),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_626),
.B(n_355),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_662),
.A2(n_365),
.B1(n_367),
.B2(n_357),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_682),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_691),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_670),
.B(n_359),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_627),
.B(n_370),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_606),
.B(n_371),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_712),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_670),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_621),
.B(n_363),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_670),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_621),
.B(n_628),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_685),
.B(n_390),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_579),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_685),
.B(n_389),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_582),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_628),
.B(n_379),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_583),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_583),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_579),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_609),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_758),
.A2(n_605),
.B(n_629),
.C(n_646),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_758),
.B(n_627),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_787),
.A2(n_652),
.B(n_648),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_781),
.B(n_659),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_717),
.A2(n_652),
.B(n_696),
.C(n_686),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_733),
.A2(n_631),
.B(n_651),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_834),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_790),
.B(n_659),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_756),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_835),
.B(n_677),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_721),
.B(n_672),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_788),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_854),
.B(n_694),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_749),
.B(n_659),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_723),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_787),
.A2(n_701),
.B(n_707),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_721),
.B(n_789),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_824),
.A2(n_644),
.B(n_609),
.Y(n_883)
);

AOI33xp33_ASAP7_75t_L g884 ( 
.A1(n_793),
.A2(n_316),
.A3(n_306),
.B1(n_364),
.B2(n_374),
.B3(n_708),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_716),
.A2(n_701),
.B(n_707),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_727),
.B(n_694),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_725),
.A2(n_686),
.B(n_306),
.C(n_374),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_739),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_742),
.B(n_604),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_856),
.A2(n_637),
.B(n_597),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_855),
.A2(n_623),
.B(n_596),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_816),
.B(n_700),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_752),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_856),
.A2(n_623),
.B(n_601),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_816),
.A2(n_589),
.B(n_596),
.C(n_656),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_727),
.B(n_708),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_742),
.B(n_610),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_846),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_825),
.B(n_622),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_SL g900 ( 
.A1(n_722),
.A2(n_601),
.B(n_637),
.C(n_584),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_752),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_825),
.A2(n_589),
.B(n_639),
.C(n_630),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_747),
.A2(n_644),
.B(n_581),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_809),
.B(n_708),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_809),
.B(n_584),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_815),
.B(n_675),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_823),
.B(n_710),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_826),
.A2(n_828),
.B(n_827),
.Y(n_908)
);

BUFx8_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_864),
.A2(n_588),
.B(n_633),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_731),
.A2(n_347),
.B(n_378),
.C(n_710),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_858),
.A2(n_812),
.B(n_821),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_811),
.A2(n_347),
.B1(n_710),
.B2(n_588),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_821),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_785),
.A2(n_633),
.B(n_710),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_823),
.B(n_633),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_815),
.B(n_675),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_842),
.A2(n_633),
.B(n_635),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_850),
.A2(n_853),
.B(n_761),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_835),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_835),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_754),
.B(n_184),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_791),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_751),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_722),
.A2(n_183),
.B(n_182),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_800),
.B(n_7),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_819),
.A2(n_178),
.B(n_160),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_734),
.A2(n_736),
.B(n_731),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_780),
.B(n_9),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_837),
.B(n_10),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_849),
.A2(n_158),
.B(n_151),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_777),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_810),
.B(n_147),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_757),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_838),
.A2(n_146),
.B(n_139),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_783),
.B(n_11),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_843),
.A2(n_127),
.B(n_116),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_760),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_767),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_851),
.A2(n_104),
.B(n_101),
.Y(n_940)
);

NOR2x1_ASAP7_75t_L g941 ( 
.A(n_738),
.B(n_743),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_724),
.B(n_12),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_833),
.A2(n_98),
.B(n_95),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_852),
.A2(n_94),
.B(n_90),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_720),
.B(n_12),
.C(n_17),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_730),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_715),
.B(n_17),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_715),
.B(n_18),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_792),
.A2(n_86),
.B(n_79),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_798),
.A2(n_77),
.B(n_70),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_718),
.B(n_19),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_803),
.B(n_66),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_813),
.A2(n_24),
.B(n_27),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_768),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_719),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_719),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_770),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_SL g958 ( 
.A(n_837),
.B(n_29),
.Y(n_958)
);

OAI321xp33_ASAP7_75t_L g959 ( 
.A1(n_729),
.A2(n_29),
.A3(n_32),
.B1(n_33),
.B2(n_35),
.C(n_36),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_814),
.A2(n_33),
.B(n_36),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_40),
.C(n_42),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_774),
.B(n_40),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_765),
.A2(n_801),
.B1(n_811),
.B2(n_775),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_741),
.Y(n_964)
);

BUFx8_ASAP7_75t_L g965 ( 
.A(n_840),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_766),
.B(n_43),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_765),
.B(n_46),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_840),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_773),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_741),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_728),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_862),
.A2(n_817),
.B(n_806),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_732),
.B(n_47),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_748),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_796),
.B(n_47),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_820),
.A2(n_52),
.B(n_53),
.Y(n_976)
);

BUFx8_ASAP7_75t_L g977 ( 
.A(n_830),
.Y(n_977)
);

NAND3xp33_ASAP7_75t_L g978 ( 
.A(n_764),
.B(n_61),
.C(n_769),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_740),
.A2(n_772),
.B1(n_726),
.B2(n_784),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_796),
.B(n_859),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_802),
.B(n_859),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_795),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_860),
.A2(n_804),
.B(n_808),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_799),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_778),
.B(n_776),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_857),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_799),
.B(n_831),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_762),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_737),
.B(n_744),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_762),
.A2(n_786),
.B(n_782),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_832),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_779),
.A2(n_750),
.B1(n_759),
.B2(n_848),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_836),
.B(n_740),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_771),
.A2(n_782),
.B(n_786),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_806),
.A2(n_817),
.B(n_745),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_772),
.B(n_841),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_753),
.A2(n_763),
.B(n_755),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_784),
.B(n_829),
.Y(n_998)
);

CKINVDCx6p67_ASAP7_75t_R g999 ( 
.A(n_818),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_797),
.B(n_845),
.C(n_822),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_844),
.B(n_805),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_735),
.A2(n_841),
.B(n_794),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_841),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_807),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_841),
.A2(n_746),
.B(n_733),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_841),
.A2(n_863),
.B(n_722),
.C(n_758),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_758),
.B(n_790),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_758),
.B(n_781),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_758),
.A2(n_725),
.B(n_717),
.C(n_721),
.Y(n_1009)
);

BUFx4f_ASAP7_75t_L g1010 ( 
.A(n_835),
.Y(n_1010)
);

OAI321xp33_ASAP7_75t_L g1011 ( 
.A1(n_758),
.A2(n_575),
.A3(n_515),
.B1(n_717),
.B2(n_721),
.C(n_479),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_758),
.B(n_781),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_742),
.A2(n_758),
.B1(n_811),
.B2(n_765),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_788),
.B(n_758),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_758),
.B(n_790),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_758),
.B(n_781),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_847),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_723),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_723),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_752),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_854),
.B(n_799),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_855),
.A2(n_716),
.B(n_787),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_788),
.B(n_758),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_861),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_1005),
.A2(n_882),
.B(n_868),
.Y(n_1025)
);

AO22x1_ASAP7_75t_L g1026 ( 
.A1(n_875),
.A2(n_973),
.B1(n_966),
.B2(n_945),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_879),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_1011),
.A2(n_1013),
.B1(n_1015),
.B2(n_1007),
.C(n_1009),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_1022),
.A2(n_994),
.B(n_990),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_880),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_1011),
.A2(n_1012),
.B(n_1016),
.C(n_1008),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1033)
);

AOI221x1_ASAP7_75t_L g1034 ( 
.A1(n_1013),
.A2(n_912),
.B1(n_896),
.B2(n_904),
.C(n_961),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_963),
.A2(n_979),
.B1(n_967),
.B2(n_993),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_1001),
.A2(n_947),
.B(n_948),
.C(n_978),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_930),
.B(n_958),
.C(n_942),
.Y(n_1037)
);

AOI221x1_ASAP7_75t_L g1038 ( 
.A1(n_912),
.A2(n_865),
.B1(n_911),
.B2(n_908),
.C(n_967),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_869),
.A2(n_998),
.B(n_889),
.C(n_897),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_979),
.A2(n_996),
.B1(n_1004),
.B2(n_866),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_983),
.A2(n_992),
.B(n_1000),
.C(n_919),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_870),
.A2(n_894),
.B(n_890),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_905),
.B(n_892),
.Y(n_1043)
);

AOI221xp5_ASAP7_75t_SL g1044 ( 
.A1(n_962),
.A2(n_936),
.B1(n_926),
.B2(n_1019),
.C(n_938),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1017),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_932),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_920),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_876),
.B(n_946),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_893),
.B(n_920),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_985),
.B(n_888),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_871),
.Y(n_1051)
);

AO31x2_ASAP7_75t_L g1052 ( 
.A1(n_895),
.A2(n_902),
.A3(n_1002),
.B(n_975),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_898),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_893),
.A2(n_878),
.B(n_867),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_924),
.B(n_934),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_939),
.B(n_954),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_957),
.B(n_969),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_885),
.A2(n_903),
.B(n_980),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_893),
.A2(n_867),
.B(n_914),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1006),
.A2(n_989),
.B(n_899),
.C(n_1018),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_898),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_SL g1062 ( 
.A1(n_949),
.A2(n_950),
.B(n_940),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_941),
.A2(n_872),
.B(n_929),
.C(n_982),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_923),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_971),
.A2(n_1021),
.B1(n_933),
.B2(n_987),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_981),
.B(n_964),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_881),
.A2(n_995),
.B(n_918),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_955),
.B(n_964),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_920),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_955),
.B(n_970),
.Y(n_1070)
);

CKINVDCx11_ASAP7_75t_R g1071 ( 
.A(n_968),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_921),
.B(n_901),
.Y(n_1072)
);

INVxp67_ASAP7_75t_SL g1073 ( 
.A(n_901),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_986),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_956),
.B(n_970),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_921),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_921),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_995),
.A2(n_1003),
.B(n_915),
.Y(n_1078)
);

BUFx8_ASAP7_75t_L g1079 ( 
.A(n_984),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_956),
.B(n_988),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1020),
.A2(n_886),
.B(n_913),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_988),
.B(n_1024),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_913),
.A2(n_927),
.B(n_931),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_SL g1084 ( 
.A1(n_975),
.A2(n_951),
.B(n_987),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_974),
.B(n_884),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_900),
.A2(n_922),
.B(n_952),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_943),
.A2(n_910),
.B(n_1021),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_935),
.A2(n_944),
.B(n_937),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1020),
.B(n_997),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1020),
.A2(n_925),
.B(n_960),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_984),
.B(n_953),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_959),
.A2(n_976),
.B(n_887),
.C(n_991),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_984),
.B(n_999),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_968),
.B(n_959),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_L g1095 ( 
.A1(n_877),
.A2(n_874),
.B(n_907),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_916),
.A2(n_907),
.B(n_877),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_916),
.A2(n_1010),
.B(n_874),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_874),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1010),
.A2(n_977),
.B(n_909),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_977),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_873),
.A2(n_882),
.B(n_1009),
.C(n_758),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_965),
.B(n_873),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_909),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_987),
.B(n_1021),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_882),
.A2(n_1009),
.B(n_1013),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_882),
.A2(n_896),
.B(n_904),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1013),
.A2(n_1012),
.B1(n_1016),
.B2(n_1008),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_882),
.B(n_758),
.C(n_721),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1011),
.A2(n_882),
.B(n_758),
.C(n_1009),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_891),
.A2(n_917),
.B(n_906),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_882),
.A2(n_758),
.B(n_721),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_882),
.A2(n_1009),
.B(n_758),
.C(n_1011),
.Y(n_1117)
);

BUFx4_ASAP7_75t_SL g1118 ( 
.A(n_874),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_901),
.Y(n_1119)
);

NAND2x1_ASAP7_75t_SL g1120 ( 
.A(n_892),
.B(n_810),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_882),
.A2(n_1009),
.B(n_758),
.C(n_1011),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_882),
.B(n_758),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_891),
.A2(n_917),
.B(n_906),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_882),
.B(n_758),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_987),
.B(n_1021),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1130)
);

AOI221x1_ASAP7_75t_L g1131 ( 
.A1(n_882),
.A2(n_758),
.B1(n_1013),
.B2(n_945),
.C(n_912),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_955),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_880),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_879),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_879),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_882),
.B(n_758),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_920),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_880),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_874),
.B(n_835),
.Y(n_1147)
);

OAI22x1_ASAP7_75t_L g1148 ( 
.A1(n_973),
.A2(n_758),
.B1(n_875),
.B2(n_1007),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_972),
.A2(n_891),
.B(n_883),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_882),
.A2(n_758),
.B(n_928),
.C(n_725),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_871),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_955),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_920),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_987),
.B(n_1021),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_920),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1031),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1140),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1053),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1122),
.A2(n_1125),
.B(n_1143),
.C(n_1115),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1107),
.A2(n_1157),
.B1(n_1150),
.B2(n_1133),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1107),
.B(n_1133),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1027),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1045),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1076),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1076),
.B(n_1047),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1137),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1112),
.B(n_1128),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1142),
.B(n_1033),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1155),
.B(n_1147),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1061),
.B(n_1137),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1139),
.B(n_1150),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1074),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_1103),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1069),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1061),
.Y(n_1179)
);

AOI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1148),
.A2(n_1113),
.B(n_1037),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1139),
.A2(n_1157),
.B1(n_1029),
.B2(n_1117),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1069),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_1071),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_1032),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1095),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_L g1186 ( 
.A(n_1121),
.B(n_1036),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1138),
.B(n_1043),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1135),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1110),
.B(n_1050),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1064),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1079),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1138),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1046),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1110),
.B(n_1050),
.Y(n_1194)
);

CKINVDCx8_ASAP7_75t_R g1195 ( 
.A(n_1103),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1145),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1103),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1048),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1147),
.B(n_1099),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1029),
.A2(n_1105),
.B1(n_1035),
.B2(n_1056),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1079),
.Y(n_1201)
);

INVx3_ASAP7_75t_SL g1202 ( 
.A(n_1100),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1105),
.A2(n_1035),
.B1(n_1055),
.B2(n_1057),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1069),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1055),
.A2(n_1056),
.B1(n_1057),
.B2(n_1094),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1038),
.A2(n_1067),
.B(n_1058),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1151),
.A2(n_1041),
.B(n_1039),
.C(n_1060),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1077),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1147),
.B(n_1098),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1120),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1152),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1026),
.B(n_1040),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1077),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1131),
.B(n_1034),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1096),
.Y(n_1216)
);

AOI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1044),
.A2(n_1091),
.B(n_1085),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1118),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1091),
.A2(n_1085),
.B1(n_1153),
.B2(n_1141),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1127),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_1049),
.B(n_1097),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1051),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1098),
.B(n_1047),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1063),
.B(n_1132),
.Y(n_1225)
);

AO22x2_ASAP7_75t_L g1226 ( 
.A1(n_1083),
.A2(n_1054),
.B1(n_1089),
.B2(n_1059),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_1098),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1077),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1066),
.B(n_1092),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1098),
.B(n_1156),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1066),
.B(n_1025),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1025),
.B(n_1082),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1068),
.A2(n_1080),
.B1(n_1070),
.B2(n_1075),
.Y(n_1233)
);

AOI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1062),
.A2(n_1089),
.B(n_1075),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1068),
.B(n_1080),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1081),
.A2(n_1049),
.B1(n_1072),
.B2(n_1088),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1154),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1088),
.A2(n_1087),
.B(n_1090),
.C(n_1086),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1154),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1119),
.B(n_1052),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1119),
.Y(n_1242)
);

INVx3_ASAP7_75t_SL g1243 ( 
.A(n_1100),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1144),
.A2(n_1156),
.B1(n_1086),
.B2(n_1154),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1072),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1144),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1102),
.B(n_1078),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1102),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1052),
.B(n_1028),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1052),
.B(n_1042),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1106),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1108),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1109),
.B(n_1124),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1084),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1114),
.B(n_1123),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1030),
.B(n_1111),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1116),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1126),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1130),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1134),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1149),
.B(n_1136),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1095),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1074),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1037),
.A2(n_882),
.B1(n_973),
.B2(n_1112),
.Y(n_1265)
);

BUFx10_ASAP7_75t_L g1266 ( 
.A(n_1074),
.Y(n_1266)
);

INVx3_ASAP7_75t_SL g1267 ( 
.A(n_1074),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1031),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1122),
.B(n_758),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1140),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1031),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1031),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1031),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1122),
.A2(n_758),
.B(n_1125),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1031),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1122),
.A2(n_1013),
.B1(n_1143),
.B2(n_1125),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1122),
.A2(n_1143),
.B1(n_1125),
.B2(n_882),
.Y(n_1283)
);

OAI321xp33_ASAP7_75t_L g1284 ( 
.A1(n_1122),
.A2(n_882),
.A3(n_758),
.B1(n_1125),
.B2(n_1143),
.C(n_1115),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1122),
.A2(n_1013),
.B1(n_1143),
.B2(n_1125),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1038),
.A2(n_1067),
.B(n_1058),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1095),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1140),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1122),
.A2(n_1143),
.B(n_1125),
.C(n_882),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1031),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1076),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1122),
.A2(n_1013),
.B1(n_1143),
.B2(n_1125),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1053),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1122),
.B(n_758),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1140),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1041),
.A2(n_1005),
.B(n_746),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1041),
.A2(n_1005),
.B(n_746),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1190),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1168),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1269),
.A2(n_1297),
.B1(n_1293),
.B2(n_1281),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1179),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1168),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1196),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1271),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1170),
.B(n_1212),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1209),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1176),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1177),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1283),
.B(n_1273),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1275),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1192),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1255),
.A2(n_1256),
.B(n_1261),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1294),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1231),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1209),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1173),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1232),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1164),
.B(n_1165),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1247),
.Y(n_1322)
);

BUFx8_ASAP7_75t_L g1323 ( 
.A(n_1168),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1250),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1240),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1292),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1193),
.Y(n_1327)
);

INVx5_ASAP7_75t_L g1328 ( 
.A(n_1222),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1283),
.A2(n_1289),
.B1(n_1175),
.B2(n_1280),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1281),
.A2(n_1293),
.B1(n_1285),
.B2(n_1265),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1203),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1183),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1247),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1203),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1188),
.Y(n_1335)
);

BUFx2_ASAP7_75t_R g1336 ( 
.A(n_1195),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1299),
.A2(n_1300),
.B(n_1260),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1292),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1252),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1222),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1249),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1173),
.B(n_1199),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1260),
.A2(n_1237),
.B(n_1216),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1215),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1189),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1285),
.A2(n_1278),
.B1(n_1186),
.B2(n_1180),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1347)
);

BUFx2_ASAP7_75t_R g1348 ( 
.A(n_1218),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1268),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1274),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1185),
.A2(n_1263),
.B(n_1287),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1279),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1226),
.A2(n_1253),
.B(n_1200),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1296),
.A2(n_1200),
.B1(n_1214),
.B2(n_1171),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1164),
.B(n_1162),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_R g1356 ( 
.A(n_1197),
.B(n_1211),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1291),
.Y(n_1357)
);

AO21x1_ASAP7_75t_L g1358 ( 
.A1(n_1181),
.A2(n_1205),
.B(n_1217),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1278),
.A2(n_1220),
.B1(n_1172),
.B2(n_1181),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1263),
.B(n_1287),
.Y(n_1360)
);

BUFx2_ASAP7_75t_R g1361 ( 
.A(n_1264),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1284),
.A2(n_1184),
.B(n_1194),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1233),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1191),
.A2(n_1267),
.B1(n_1201),
.B2(n_1243),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1174),
.B(n_1205),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1207),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1226),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1198),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1160),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1234),
.A2(n_1259),
.B(n_1229),
.Y(n_1370)
);

INVx4_ASAP7_75t_SL g1371 ( 
.A(n_1222),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1235),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1251),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1206),
.A2(n_1286),
.B(n_1225),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1206),
.A2(n_1286),
.B(n_1219),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1245),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1251),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1159),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1187),
.A2(n_1248),
.B1(n_1210),
.B2(n_1254),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1221),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1284),
.A2(n_1210),
.B1(n_1202),
.B2(n_1223),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1253),
.A2(n_1257),
.B(n_1236),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1199),
.A2(n_1270),
.B1(n_1298),
.B2(n_1288),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1266),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1292),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1245),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1242),
.Y(n_1387)
);

BUFx8_ASAP7_75t_SL g1388 ( 
.A(n_1166),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1259),
.B(n_1244),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1246),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1224),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1266),
.A2(n_1161),
.B1(n_1163),
.B2(n_1290),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1167),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1161),
.A2(n_1163),
.B1(n_1290),
.B2(n_1282),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1258),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1258),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1272),
.A2(n_1295),
.B1(n_1282),
.B2(n_1199),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1272),
.A2(n_1295),
.B1(n_1227),
.B2(n_1230),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1245),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1240),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1240),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1262),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1244),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1239),
.A2(n_1169),
.B(n_1230),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1246),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1246),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1182),
.A2(n_1238),
.B1(n_1178),
.B2(n_1213),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1178),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1213),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1204),
.A2(n_1208),
.B(n_1228),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1177),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1192),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1247),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1269),
.A2(n_875),
.B1(n_882),
.B2(n_758),
.Y(n_1414)
);

AO21x1_ASAP7_75t_L g1415 ( 
.A1(n_1186),
.A2(n_1113),
.B(n_882),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1241),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1179),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1283),
.A2(n_882),
.B1(n_958),
.B2(n_930),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1158),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1190),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1170),
.B(n_1212),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1186),
.A2(n_1113),
.B(n_882),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1190),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1283),
.A2(n_1122),
.B1(n_1143),
.B2(n_1125),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1269),
.A2(n_882),
.B1(n_1037),
.B2(n_973),
.Y(n_1425)
);

AO21x1_ASAP7_75t_L g1426 ( 
.A1(n_1186),
.A2(n_1113),
.B(n_882),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1269),
.A2(n_958),
.B1(n_930),
.B2(n_758),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1240),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1190),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1241),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1310),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1339),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1324),
.B(n_1321),
.Y(n_1433)
);

AO21x1_ASAP7_75t_L g1434 ( 
.A1(n_1418),
.A2(n_1362),
.B(n_1381),
.Y(n_1434)
);

BUFx4f_ASAP7_75t_SL g1435 ( 
.A(n_1332),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1324),
.B(n_1321),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1365),
.B(n_1355),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1412),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1347),
.B(n_1312),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1374),
.A2(n_1375),
.B(n_1358),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1328),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1358),
.A2(n_1367),
.B(n_1337),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1416),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1329),
.B(n_1424),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1416),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1365),
.B(n_1355),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1412),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1317),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1414),
.B(n_1354),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1317),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1368),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1344),
.B(n_1430),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1344),
.B(n_1331),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1304),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1367),
.A2(n_1353),
.B(n_1363),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1389),
.B(n_1340),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1369),
.B(n_1310),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1343),
.A2(n_1315),
.B(n_1351),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1308),
.B(n_1421),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1382),
.A2(n_1315),
.B(n_1353),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1331),
.A2(n_1334),
.B(n_1343),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1320),
.Y(n_1463)
);

INVx8_ASAP7_75t_L g1464 ( 
.A(n_1401),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1351),
.A2(n_1404),
.B(n_1389),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1341),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1327),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1415),
.A2(n_1422),
.B(n_1426),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1427),
.A2(n_1425),
.B1(n_1303),
.B2(n_1330),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1341),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1322),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1403),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1403),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1360),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1322),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1415),
.A2(n_1422),
.B(n_1426),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1345),
.A2(n_1346),
.B(n_1377),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1333),
.B(n_1413),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1373),
.A2(n_1377),
.B(n_1402),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1333),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1371),
.B(n_1413),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1413),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1393),
.B(n_1316),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1340),
.B(n_1370),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1417),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1370),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1345),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1378),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1373),
.A2(n_1359),
.B(n_1366),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1336),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1340),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1335),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1342),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1352),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1342),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1371),
.B(n_1342),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1371),
.B(n_1395),
.Y(n_1497)
);

INVxp33_ASAP7_75t_L g1498 ( 
.A(n_1388),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1371),
.B(n_1396),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1349),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1372),
.B(n_1306),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1350),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1383),
.A2(n_1357),
.B(n_1387),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1306),
.B(n_1419),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1379),
.A2(n_1392),
.B(n_1307),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1309),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1301),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1444),
.A2(n_1319),
.B1(n_1318),
.B2(n_1309),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1438),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1460),
.B(n_1313),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1447),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1432),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1437),
.B(n_1380),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1437),
.B(n_1319),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1439),
.B(n_1318),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1431),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1451),
.B(n_1318),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1446),
.B(n_1319),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1456),
.B(n_1319),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1452),
.B(n_1318),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1457),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1481),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1446),
.B(n_1319),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1481),
.B(n_1496),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1469),
.A2(n_1397),
.B1(n_1394),
.B2(n_1398),
.C(n_1301),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1456),
.B(n_1309),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1486),
.A2(n_1459),
.B(n_1461),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1449),
.A2(n_1384),
.B1(n_1361),
.B2(n_1420),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1456),
.B(n_1429),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1456),
.B(n_1429),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1435),
.B(n_1420),
.Y(n_1536)
);

BUFx2_ASAP7_75t_R g1537 ( 
.A(n_1506),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1466),
.B(n_1386),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1479),
.B(n_1408),
.Y(n_1542)
);

AND2x4_ASAP7_75t_SL g1543 ( 
.A(n_1496),
.B(n_1391),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1479),
.B(n_1408),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1505),
.A2(n_1410),
.B(n_1384),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1485),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1466),
.B(n_1470),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_R g1548 ( 
.A(n_1431),
.B(n_1332),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1488),
.B(n_1386),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1399),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1486),
.B(n_1409),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1462),
.B(n_1409),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1464),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1434),
.A2(n_1364),
.B1(n_1311),
.B2(n_1305),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1457),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1501),
.B(n_1376),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1462),
.B(n_1410),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1471),
.B(n_1376),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1442),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1545),
.B(n_1483),
.C(n_1467),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1535),
.B(n_1434),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1554),
.A2(n_1490),
.B1(n_1507),
.B2(n_1457),
.C(n_1478),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1492),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1546),
.B(n_1494),
.Y(n_1564)
);

NOR3xp33_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1458),
.C(n_1491),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1482),
.C(n_1480),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1527),
.A2(n_1498),
.B(n_1496),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1475),
.C(n_1473),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1516),
.A2(n_1311),
.B1(n_1457),
.B2(n_1477),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1509),
.A2(n_1468),
.B1(n_1476),
.B2(n_1489),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1534),
.C(n_1538),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1511),
.B(n_1448),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1533),
.B(n_1475),
.C(n_1473),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1472),
.C(n_1487),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1535),
.A2(n_1474),
.B(n_1465),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1510),
.B(n_1450),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_1442),
.Y(n_1578)
);

NOR3xp33_ASAP7_75t_L g1579 ( 
.A(n_1515),
.B(n_1491),
.C(n_1356),
.Y(n_1579)
);

AND2x4_ASAP7_75t_SL g1580 ( 
.A(n_1526),
.B(n_1497),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1538),
.A2(n_1478),
.B1(n_1487),
.B2(n_1407),
.C(n_1500),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1547),
.B(n_1442),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1539),
.B(n_1472),
.C(n_1477),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1442),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_L g1585 ( 
.A(n_1539),
.B(n_1491),
.C(n_1325),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1508),
.A2(n_1493),
.B1(n_1495),
.B2(n_1499),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1517),
.B(n_1502),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1463),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1512),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1537),
.A2(n_1493),
.B1(n_1495),
.B2(n_1497),
.Y(n_1590)
);

NOR3xp33_ASAP7_75t_L g1591 ( 
.A(n_1522),
.B(n_1491),
.C(n_1325),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1536),
.A2(n_1302),
.B1(n_1305),
.B2(n_1385),
.C(n_1326),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1428),
.C(n_1504),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1516),
.A2(n_1495),
.B1(n_1499),
.B2(n_1497),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1512),
.Y(n_1596)
);

NAND2xp33_ASAP7_75t_SL g1597 ( 
.A(n_1548),
.B(n_1441),
.Y(n_1597)
);

OAI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1519),
.A2(n_1529),
.B(n_1513),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1513),
.B(n_1453),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1443),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1543),
.A2(n_1497),
.B(n_1499),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1521),
.B(n_1462),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1541),
.B(n_1443),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1604)
);

OAI21xp33_ASAP7_75t_L g1605 ( 
.A1(n_1519),
.A2(n_1454),
.B(n_1445),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1521),
.B(n_1462),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1559),
.B(n_1523),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1578),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1571),
.B(n_1552),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1589),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1580),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1582),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1584),
.B(n_1530),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1575),
.B(n_1524),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1602),
.B(n_1530),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1530),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1606),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1606),
.B(n_1530),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1604),
.B(n_1598),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1572),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1577),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1561),
.B(n_1441),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1583),
.B(n_1603),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1529),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_1542),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1561),
.A2(n_1476),
.B1(n_1468),
.B2(n_1489),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1573),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1570),
.B(n_1440),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1570),
.B(n_1440),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1580),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1588),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1566),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1587),
.B(n_1542),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1544),
.Y(n_1641)
);

INVxp33_ASAP7_75t_L g1642 ( 
.A(n_1565),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1597),
.B(n_1526),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1642),
.B(n_1567),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1611),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1611),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1614),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1629),
.B(n_1563),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1614),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1639),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1608),
.B(n_1524),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_SL g1655 ( 
.A(n_1643),
.B(n_1601),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1524),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1639),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1624),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1624),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1627),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1624),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1638),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1616),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1640),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1564),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1608),
.B(n_1585),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1612),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1638),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1629),
.B(n_1599),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1638),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1609),
.B(n_1551),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1607),
.B(n_1558),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1618),
.B(n_1593),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1642),
.B(n_1592),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1607),
.B(n_1558),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1616),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1609),
.B(n_1551),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1615),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1609),
.B(n_1605),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1610),
.B(n_1525),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1640),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1610),
.B(n_1525),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1610),
.B(n_1637),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1643),
.B(n_1597),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1637),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1655),
.B(n_1681),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1645),
.Y(n_1691)
);

OAI211xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1677),
.A2(n_1626),
.B(n_1633),
.C(n_1635),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1633),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1644),
.B(n_1633),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

OR4x1_ASAP7_75t_L g1696 ( 
.A(n_1667),
.B(n_1626),
.C(n_1581),
.D(n_1562),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1626),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1646),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1646),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1665),
.B(n_1641),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1648),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1650),
.B(n_1631),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1648),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1641),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1688),
.B(n_1631),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1667),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1649),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1681),
.A2(n_1569),
.B1(n_1586),
.B2(n_1618),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1649),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1666),
.B(n_1630),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1651),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1676),
.B(n_1618),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1676),
.B(n_1618),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1685),
.B(n_1630),
.Y(n_1717)
);

NAND2x2_ASAP7_75t_L g1718 ( 
.A(n_1683),
.B(n_1411),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1669),
.B(n_1613),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1647),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1651),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1654),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1654),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1670),
.B(n_1630),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1666),
.B(n_1623),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1618),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1658),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1676),
.A2(n_1635),
.B(n_1627),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1669),
.A2(n_1618),
.B1(n_1590),
.B2(n_1636),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1687),
.B(n_1612),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1670),
.B(n_1684),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1683),
.B(n_1625),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1647),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1690),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1689),
.B(n_1687),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1732),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1691),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1653),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1695),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1698),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1712),
.B(n_1653),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1699),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1701),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1702),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1694),
.A2(n_1660),
.B(n_1627),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1704),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1706),
.B(n_1686),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1720),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1731),
.B(n_1674),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1692),
.A2(n_1718),
.B1(n_1706),
.B2(n_1709),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1720),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1713),
.B(n_1656),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1715),
.B(n_1656),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1708),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1692),
.A2(n_1636),
.B1(n_1634),
.B2(n_1627),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1700),
.B(n_1684),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1697),
.B(n_1674),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1710),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1675),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1714),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1724),
.B(n_1680),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1766)
);

AND2x4_ASAP7_75t_SL g1767 ( 
.A(n_1715),
.B(n_1632),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1703),
.B(n_1680),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1659),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1721),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1733),
.B(n_1678),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1753),
.A2(n_1718),
.B1(n_1729),
.B2(n_1632),
.Y(n_1773)
);

XNOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1735),
.B(n_1696),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1767),
.A2(n_1696),
.B1(n_1733),
.B2(n_1627),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1763),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1742),
.B(n_1705),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1769),
.B(n_1727),
.C(n_1730),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1769),
.A2(n_1716),
.B1(n_1726),
.B2(n_1636),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1759),
.A2(n_1726),
.B(n_1716),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1745),
.Y(n_1782)
);

AOI32xp33_ASAP7_75t_L g1783 ( 
.A1(n_1767),
.A2(n_1716),
.A3(n_1726),
.B1(n_1634),
.B2(n_1717),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1738),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1737),
.A2(n_1612),
.B1(n_1348),
.B2(n_1722),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1738),
.Y(n_1787)
);

AOI31xp33_ASAP7_75t_L g1788 ( 
.A1(n_1752),
.A2(n_1594),
.A3(n_1723),
.B(n_1634),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1760),
.B(n_1659),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1740),
.B(n_1661),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1737),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1734),
.C(n_1661),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1740),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1741),
.B(n_1744),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1741),
.B(n_1682),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1678),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1747),
.A2(n_1668),
.B(n_1662),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1763),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1744),
.Y(n_1799)
);

AOI322xp5_ASAP7_75t_L g1800 ( 
.A1(n_1749),
.A2(n_1622),
.A3(n_1620),
.B1(n_1619),
.B2(n_1617),
.C1(n_1621),
.C2(n_1623),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1791),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1782),
.B(n_1772),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1794),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1776),
.B(n_1779),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1775),
.B(n_1739),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1777),
.B(n_1739),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1774),
.B(n_1743),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1776),
.B(n_1761),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.B(n_1761),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1794),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1798),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1796),
.B(n_1743),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1785),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1792),
.B(n_1746),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1786),
.B(n_1768),
.Y(n_1815)
);

CKINVDCx16_ASAP7_75t_R g1816 ( 
.A(n_1773),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1787),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1784),
.A2(n_1751),
.B1(n_1767),
.B2(n_1765),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1793),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1778),
.B(n_1757),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1757),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1799),
.B(n_1766),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1801),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1816),
.A2(n_1781),
.B1(n_1748),
.B2(n_1758),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1804),
.A2(n_1783),
.B1(n_1788),
.B2(n_1797),
.C(n_1789),
.Y(n_1825)
);

AOI211xp5_ASAP7_75t_L g1826 ( 
.A1(n_1815),
.A2(n_1762),
.B(n_1746),
.C(n_1758),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1808),
.A2(n_1807),
.B1(n_1818),
.B2(n_1802),
.C(n_1801),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1803),
.A2(n_1810),
.B1(n_1820),
.B2(n_1811),
.C(n_1822),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1814),
.A2(n_1768),
.B1(n_1751),
.B2(n_1765),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1809),
.A2(n_1800),
.B1(n_1790),
.B2(n_1764),
.C(n_1771),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1809),
.B(n_1755),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1821),
.A2(n_1790),
.B(n_1795),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1811),
.B(n_1795),
.C(n_1762),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1820),
.B(n_1755),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1805),
.B(n_1748),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1821),
.A2(n_1771),
.B(n_1764),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_SL g1837 ( 
.A(n_1826),
.B(n_1805),
.C(n_1806),
.D(n_1812),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_L g1838 ( 
.A(n_1827),
.B(n_1813),
.C(n_1810),
.Y(n_1838)
);

NOR3xp33_ASAP7_75t_L g1839 ( 
.A(n_1829),
.B(n_1803),
.C(n_1817),
.Y(n_1839)
);

NAND4xp75_ASAP7_75t_L g1840 ( 
.A(n_1828),
.B(n_1823),
.C(n_1824),
.D(n_1831),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1834),
.B(n_1806),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1835),
.B(n_1812),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1825),
.B(n_1819),
.C(n_1817),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1830),
.A2(n_1819),
.B1(n_1621),
.B2(n_1612),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1833),
.Y(n_1845)
);

NOR3x1_ASAP7_75t_L g1846 ( 
.A(n_1836),
.B(n_1682),
.C(n_1668),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1832),
.A2(n_1770),
.B(n_1754),
.C(n_1750),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1840),
.B(n_1754),
.C(n_1750),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1839),
.B(n_1754),
.C(n_1750),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1842),
.B(n_1770),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1837),
.B(n_1323),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1841),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1845),
.B(n_1844),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1850),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1849),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1852),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_SL g1857 ( 
.A(n_1851),
.B(n_1838),
.C(n_1843),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1848),
.Y(n_1858)
);

OR2x6_ASAP7_75t_L g1859 ( 
.A(n_1853),
.B(n_1411),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1851),
.A2(n_1847),
.B1(n_1770),
.B2(n_1846),
.Y(n_1860)
);

NOR3xp33_ASAP7_75t_L g1861 ( 
.A(n_1857),
.B(n_1326),
.C(n_1302),
.Y(n_1861)
);

INVx3_ASAP7_75t_SL g1862 ( 
.A(n_1859),
.Y(n_1862)
);

OAI211xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1858),
.A2(n_1855),
.B(n_1854),
.C(n_1856),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1860),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1857),
.A2(n_1671),
.B(n_1662),
.Y(n_1865)
);

NOR2xp67_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1428),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1862),
.B(n_1647),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1863),
.B(n_1663),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1866),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1864),
.A2(n_1679),
.B1(n_1663),
.B2(n_1671),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1867),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1869),
.B(n_1861),
.Y(n_1872)
);

NOR4xp25_ASAP7_75t_SL g1873 ( 
.A(n_1871),
.B(n_1868),
.C(n_1865),
.D(n_1870),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1873),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1873),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1875),
.B(n_1872),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1874),
.B(n_1872),
.Y(n_1877)
);

OR2x6_ASAP7_75t_L g1878 ( 
.A(n_1876),
.B(n_1877),
.Y(n_1878)
);

AOI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_1400),
.B(n_1663),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_1323),
.B1(n_1390),
.B2(n_1338),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1672),
.B1(n_1338),
.B2(n_1385),
.C(n_1679),
.Y(n_1881)
);

AOI211xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1401),
.B(n_1405),
.C(n_1406),
.Y(n_1882)
);


endmodule