module fake_jpeg_3292_n_498 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_498);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_498;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_49),
.B(n_48),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_54),
.Y(n_105)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_0),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_82),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_40),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_84),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_1),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_20),
.B(n_1),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_R g91 ( 
.A(n_40),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_42),
.Y(n_132)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_43),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_47),
.B1(n_27),
.B2(n_45),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_97),
.A2(n_134),
.B1(n_88),
.B2(n_5),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_46),
.B1(n_18),
.B2(n_29),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_99),
.A2(n_133),
.B1(n_4),
.B2(n_5),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_47),
.C(n_38),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_100),
.B(n_6),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_47),
.B1(n_31),
.B2(n_46),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_104),
.A2(n_136),
.B1(n_147),
.B2(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_28),
.B1(n_45),
.B2(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_119),
.A2(n_125),
.B1(n_148),
.B2(n_7),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_28),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_48),
.B1(n_43),
.B2(n_20),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_53),
.A2(n_29),
.B1(n_42),
.B2(n_18),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_68),
.A2(n_93),
.B1(n_89),
.B2(n_65),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_70),
.A2(n_31),
.B1(n_42),
.B2(n_29),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_51),
.A2(n_19),
.B(n_42),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_84),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_31),
.B1(n_42),
.B2(n_29),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_56),
.A2(n_24),
.B1(n_37),
.B2(n_19),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_37),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_154),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_94),
.A2(n_29),
.B1(n_24),
.B2(n_19),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_79),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_156),
.Y(n_255)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_105),
.B(n_58),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_161),
.B(n_166),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

OR2x2_ASAP7_75t_SL g163 ( 
.A(n_100),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_163),
.Y(n_230)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_165),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_62),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_62),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_170),
.Y(n_228)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_74),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_76),
.B1(n_83),
.B2(n_80),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_171),
.A2(n_173),
.B1(n_205),
.B2(n_145),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_77),
.B1(n_73),
.B2(n_72),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_67),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_63),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_130),
.B(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_180),
.B(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_185),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_4),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_190),
.Y(n_247)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_191),
.A2(n_211),
.B(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_127),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_192),
.B(n_201),
.Y(n_262)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_15),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_106),
.B(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_201),
.B(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_99),
.A2(n_133),
.B1(n_102),
.B2(n_109),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_203),
.B1(n_113),
.B2(n_108),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_102),
.B(n_7),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_143),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_134),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g204 ( 
.A(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_103),
.A2(n_109),
.B1(n_150),
.B2(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_206),
.B(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_121),
.B(n_7),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_113),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_97),
.B1(n_119),
.B2(n_129),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_219),
.B1(n_233),
.B2(n_234),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_217),
.A2(n_218),
.B(n_231),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_199),
.B1(n_198),
.B2(n_211),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_129),
.B1(n_141),
.B2(n_101),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_221),
.B(n_262),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_138),
.B1(n_143),
.B2(n_150),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_232),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_163),
.A2(n_141),
.B1(n_101),
.B2(n_145),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_164),
.A2(n_108),
.B1(n_135),
.B2(n_140),
.Y(n_234)
);

NAND2x1p5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_236),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_170),
.A2(n_137),
.B1(n_135),
.B2(n_138),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_238),
.A2(n_245),
.B1(n_249),
.B2(n_253),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_158),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_193),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_204),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_137),
.B1(n_114),
.B2(n_12),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_190),
.A2(n_186),
.B1(n_167),
.B2(n_162),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_190),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_253),
.B1(n_216),
.B2(n_244),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_169),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_297),
.C(n_258),
.Y(n_308)
);

AOI22x1_ASAP7_75t_SL g264 ( 
.A1(n_249),
.A2(n_186),
.B1(n_206),
.B2(n_212),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_271),
.B1(n_282),
.B2(n_288),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_186),
.B1(n_189),
.B2(n_210),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_265),
.A2(n_270),
.B1(n_276),
.B2(n_283),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_175),
.B(n_174),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_267),
.A2(n_299),
.B(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_273),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_157),
.B1(n_177),
.B2(n_165),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_184),
.B1(n_187),
.B2(n_156),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_256),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_222),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_274),
.A2(n_279),
.B(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_218),
.A2(n_168),
.B1(n_183),
.B2(n_159),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_204),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_277),
.A2(n_278),
.B(n_280),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_208),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_233),
.B(n_13),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_14),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_14),
.B1(n_228),
.B2(n_217),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_240),
.A2(n_14),
.B1(n_228),
.B2(n_236),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_229),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_284),
.B(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_221),
.B(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_236),
.B(n_257),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_227),
.B(n_252),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_290),
.B(n_301),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_248),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_238),
.A2(n_248),
.B1(n_219),
.B2(n_245),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_293),
.A2(n_273),
.B1(n_295),
.B2(n_292),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_227),
.A2(n_261),
.B(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_225),
.B1(n_261),
.B2(n_215),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_255),
.B(n_241),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_225),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_251),
.B(n_214),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_300),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_237),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_234),
.A2(n_223),
.B1(n_254),
.B2(n_214),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_306),
.B1(n_307),
.B2(n_224),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_242),
.A2(n_258),
.B(n_241),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_223),
.A2(n_254),
.B1(n_235),
.B2(n_260),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_235),
.A2(n_260),
.B1(n_256),
.B2(n_242),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_308),
.B(n_309),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_313),
.B(n_347),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_255),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_317),
.C(n_331),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_250),
.C(n_224),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_299),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_324),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_265),
.B1(n_279),
.B2(n_282),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_285),
.A2(n_266),
.B1(n_305),
.B2(n_293),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_336),
.B1(n_338),
.B2(n_303),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_276),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_297),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_339),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_289),
.C(n_263),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_267),
.B(n_294),
.C(n_269),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_341),
.C(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_266),
.B1(n_305),
.B2(n_279),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_279),
.B1(n_288),
.B2(n_264),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_296),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_290),
.B(n_302),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_302),
.C(n_278),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_346),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_274),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_341),
.C(n_308),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_287),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_296),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_348),
.B(n_380),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_337),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_356),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_361),
.B1(n_367),
.B2(n_324),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_369),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_330),
.B(n_270),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_304),
.B(n_281),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_359),
.B(n_351),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_362),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_306),
.B(n_300),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_300),
.B1(n_336),
.B2(n_338),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_323),
.B(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_339),
.B1(n_346),
.B2(n_347),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_309),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_373),
.C(n_317),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_311),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_311),
.B(n_344),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_345),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_383),
.B1(n_392),
.B2(n_402),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_352),
.A2(n_324),
.B1(n_313),
.B2(n_340),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_371),
.C(n_350),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_389),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_333),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_340),
.B1(n_315),
.B2(n_329),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_315),
.B1(n_322),
.B2(n_329),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_399),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_362),
.B(n_332),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_395),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_348),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_379),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_350),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_377),
.A2(n_375),
.B1(n_355),
.B2(n_354),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_363),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_400),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_363),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_372),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_367),
.A2(n_354),
.B1(n_351),
.B2(n_365),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_404),
.B(n_359),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_349),
.A2(n_366),
.B1(n_355),
.B2(n_356),
.Y(n_404)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_403),
.B(n_383),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_431),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_404),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_413),
.B(n_388),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_430),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_398),
.C(n_389),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_418),
.C(n_423),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_405),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_370),
.C(n_373),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_391),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_422),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_391),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_370),
.C(n_357),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_424),
.Y(n_439)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_425),
.Y(n_443)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_429),
.Y(n_449)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_360),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_364),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_432),
.A2(n_410),
.B(n_427),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_444),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_416),
.B(n_388),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_437),
.Y(n_460)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_419),
.B(n_397),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_421),
.A2(n_393),
.B1(n_382),
.B2(n_405),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_440),
.A2(n_442),
.B1(n_431),
.B2(n_425),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_392),
.B1(n_408),
.B2(n_385),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_397),
.Y(n_444)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_396),
.A3(n_406),
.B1(n_407),
.B2(n_376),
.C1(n_378),
.C2(n_374),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_448),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_396),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_406),
.C(n_407),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_450),
.B(n_430),
.C(n_423),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_452),
.B(n_455),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_415),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_457),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_447),
.C(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_417),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_456),
.B(n_458),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_412),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_420),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_432),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_465),
.C(n_409),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_424),
.B(n_427),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_464),
.B1(n_443),
.B2(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_412),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_450),
.C(n_447),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_467),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_449),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_440),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_468),
.B(n_454),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_470),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_436),
.B1(n_442),
.B2(n_445),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_472),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_459),
.A2(n_409),
.B(n_426),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_463),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_473),
.B(n_452),
.CI(n_462),
.CON(n_479),
.SN(n_479)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_476),
.B(n_451),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_482),
.B(n_474),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_453),
.C(n_465),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_484),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_489),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_481),
.A2(n_475),
.B(n_471),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_486),
.A2(n_477),
.B(n_484),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_464),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_491),
.A2(n_479),
.B(n_487),
.C(n_490),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_483),
.C(n_477),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_492),
.Y(n_494)
);

MAJx2_ASAP7_75t_L g495 ( 
.A(n_493),
.B(n_457),
.C(n_461),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_494),
.C(n_472),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_428),
.Y(n_498)
);


endmodule