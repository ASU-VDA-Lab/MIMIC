module fake_jpeg_6736_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_19),
.CON(n_50),
.SN(n_50)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_35),
.B1(n_20),
.B2(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_35),
.B1(n_20),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_63),
.B1(n_20),
.B2(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_35),
.B1(n_20),
.B2(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_28),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_74),
.C(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_76),
.B(n_79),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_62),
.B(n_24),
.Y(n_116)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_38),
.B1(n_37),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_83),
.B1(n_59),
.B2(n_61),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_85),
.Y(n_119)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_99),
.B1(n_59),
.B2(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_93),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_97),
.Y(n_127)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_68),
.C(n_49),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_106),
.C(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_107),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_25),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_115),
.B(n_34),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_34),
.Y(n_148)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_69),
.C(n_63),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_60),
.B(n_53),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_64),
.B1(n_82),
.B2(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_114),
.B1(n_122),
.B2(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_42),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_72),
.C(n_29),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_64),
.B1(n_66),
.B2(n_82),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_142),
.B1(n_144),
.B2(n_66),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_134),
.B1(n_137),
.B2(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_145),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_78),
.B1(n_84),
.B2(n_86),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_91),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_26),
.B(n_31),
.Y(n_165)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_72),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_138),
.B(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_86),
.B1(n_51),
.B2(n_52),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_23),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_99),
.B1(n_88),
.B2(n_93),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_88),
.B1(n_85),
.B2(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_24),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.C(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_152),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_72),
.C(n_45),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_23),
.B(n_25),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_120),
.B(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_72),
.B(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_104),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_173),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_145),
.B(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_177),
.C(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_128),
.B1(n_127),
.B2(n_111),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_166),
.B1(n_176),
.B2(n_156),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_138),
.B(n_121),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_43),
.B1(n_29),
.B2(n_24),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_138),
.B1(n_129),
.B2(n_125),
.Y(n_212)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_29),
.B1(n_124),
.B2(n_113),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_109),
.C(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_17),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_17),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_156),
.C(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_102),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_155),
.A3(n_151),
.B1(n_132),
.B2(n_142),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_158),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_137),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_214),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_197),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_203),
.B(n_207),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_131),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_208),
.C(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_150),
.B1(n_155),
.B2(n_152),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_212),
.B1(n_160),
.B2(n_180),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_209),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_154),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_170),
.B1(n_181),
.B2(n_172),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_218),
.B1(n_222),
.B2(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_210),
.B1(n_193),
.B2(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_233),
.C(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_164),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_229),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_226),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_232),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_172),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_175),
.B(n_161),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_238),
.B(n_240),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_158),
.C(n_173),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_235),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_173),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_166),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_189),
.A2(n_178),
.B(n_171),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_17),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_187),
.B1(n_188),
.B2(n_207),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_217),
.B(n_225),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_199),
.C(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_267)
);

OAI22x1_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_200),
.B1(n_198),
.B2(n_209),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_2),
.B(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_191),
.C(n_179),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_191),
.C(n_183),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_129),
.B1(n_108),
.B2(n_102),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_262),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_129),
.C(n_139),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.C(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_139),
.C(n_121),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_227),
.C(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_231),
.B1(n_241),
.B2(n_32),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_21),
.B1(n_32),
.B2(n_22),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_21),
.B1(n_32),
.B2(n_22),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_22),
.B1(n_9),
.B2(n_10),
.Y(n_281)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_247),
.C(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_284),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_9),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_0),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_275),
.B(n_5),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_282),
.B1(n_10),
.B2(n_14),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_287),
.C(n_291),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_246),
.C(n_247),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_245),
.B1(n_254),
.B2(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_257),
.C(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_10),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_283),
.B(n_13),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_295),
.Y(n_308)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_9),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_269),
.B1(n_283),
.B2(n_273),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_273),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_280),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_311),
.B(n_313),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_270),
.B1(n_268),
.B2(n_12),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_16),
.B1(n_8),
.B2(n_11),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_4),
.C(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_294),
.C(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_4),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_12),
.B(n_14),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_324),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_321),
.B(n_311),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_295),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_6),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_308),
.A2(n_286),
.B(n_297),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_285),
.C(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_312),
.C(n_305),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_301),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_327),
.B(n_317),
.Y(n_337)
);

OA21x2_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_309),
.B(n_8),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_329),
.B(n_330),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_11),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_13),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_16),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_327),
.B(n_316),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_328),
.C(n_320),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_337),
.C(n_319),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_333),
.B(n_336),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_339),
.B(n_332),
.C(n_331),
.D(n_7),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_6),
.B(n_7),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);


endmodule