module fake_jpeg_17867_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_20),
.Y(n_24)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_6),
.B(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_21),
.B1(n_8),
.B2(n_11),
.Y(n_27)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_4),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_10),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_20),
.B(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_19),
.B1(n_15),
.B2(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_19),
.B(n_8),
.C(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_34),
.B1(n_15),
.B2(n_22),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_24),
.B(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_11),
.C(n_13),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_34),
.C(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_11),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_38),
.B(n_32),
.Y(n_44)
);

AO221x1_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B1(n_43),
.B2(n_35),
.C(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_13),
.Y(n_46)
);


endmodule