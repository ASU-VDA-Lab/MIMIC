module fake_jpeg_31421_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_8),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_46),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_40),
.B(n_18),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_28),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_18),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_24),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_41),
.B1(n_34),
.B2(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_42),
.B1(n_15),
.B2(n_17),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_77),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_60),
.B1(n_53),
.B2(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_74),
.B1(n_62),
.B2(n_56),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_27),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_27),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_68),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_66),
.C(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_74),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_74),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_47),
.B(n_26),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_103),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_79),
.B1(n_51),
.B2(n_67),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_85),
.B1(n_73),
.B2(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_111),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_95),
.C(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_103),
.C(n_87),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_101),
.C(n_98),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_93),
.C(n_85),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_112),
.C(n_93),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_105),
.B1(n_110),
.B2(n_113),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_112),
.B1(n_54),
.B2(n_50),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_128),
.Y(n_130)
);

AOI31xp67_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_112),
.A3(n_26),
.B(n_10),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_120),
.C(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_54),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_7),
.B(n_11),
.C(n_4),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_7),
.B(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_4),
.Y(n_135)
);


endmodule