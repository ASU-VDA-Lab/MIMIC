module real_jpeg_14841_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_46),
.B1(n_64),
.B2(n_66),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_27),
.C(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_28),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_4),
.B(n_51),
.C(n_54),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_61),
.C(n_66),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_19),
.B1(n_20),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_35),
.B1(n_64),
.B2(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_14),
.B(n_263),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_10),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_22),
.B1(n_54),
.B2(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_22),
.B1(n_64),
.B2(n_66),
.Y(n_88)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_38),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_37),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_32),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_32),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_23),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_20),
.B(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_30),
.B(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_32),
.B(n_40),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_45),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_72),
.B(n_262),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_70),
.C(n_71),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_41),
.A2(n_42),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_57),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_44),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_43),
.B(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_43),
.A2(n_44),
.B1(n_93),
.B2(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_43),
.A2(n_44),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI211xp5_ASAP7_75t_SL g162 ( 
.A1(n_43),
.A2(n_89),
.B(n_110),
.C(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_43),
.A2(n_44),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_43),
.A2(n_93),
.B(n_117),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_43),
.A2(n_44),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_43),
.A2(n_44),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_44),
.B(n_81),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_44),
.B(n_58),
.C(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_44),
.B(n_247),
.C(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_46),
.B(n_101),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_46),
.B(n_87),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_47),
.A2(n_57),
.B1(n_58),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_47),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_82),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_53),
.B(n_56),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_53),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_53),
.Y(n_198)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_54),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_57),
.A2(n_58),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_69),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_67),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_68),
.Y(n_67)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_67),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_67),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_64),
.B(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_70),
.B(n_71),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_256),
.B(n_261),
.Y(n_72)
);

AOI21x1_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_230),
.B(n_253),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_128),
.B(n_229),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_111),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_76),
.B(n_111),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_92),
.C(n_103),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_91),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_78),
.A2(n_79),
.B1(n_105),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_78),
.A2(n_79),
.B1(n_142),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_138),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_146),
.C(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_80),
.A2(n_81),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_81),
.B(n_138),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_81),
.A2(n_138),
.B(n_175),
.C(n_180),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_104),
.B(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_89),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_89),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_89),
.A2(n_106),
.B1(n_138),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_89),
.A2(n_138),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_89),
.A2(n_138),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_89),
.A2(n_138),
.B1(n_192),
.B2(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_89),
.B(n_146),
.C(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_89),
.B(n_182),
.C(n_186),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_102),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_97),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_109),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_109),
.B(n_142),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_127),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_116),
.B(n_121),
.C(n_127),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_126),
.A2(n_234),
.B1(n_235),
.B2(n_240),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_148),
.B(n_228),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_130),
.B(n_132),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_140),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_140),
.A2(n_141),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_147),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_147),
.B1(n_157),
.B2(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_147),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_146),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_146),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_147),
.B(n_208),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_169),
.B(n_222),
.C(n_227),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_153),
.B1(n_175),
.B2(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_216),
.B(n_221),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_188),
.B(n_215),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_211),
.B(n_214),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_200),
.B(n_210),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_242),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_242),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_241),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_240),
.C(n_241),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_252),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_260),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);


endmodule