module real_jpeg_5645_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_1),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_1),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_1),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_1),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_1),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_2),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_3),
.B(n_85),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_5),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_5),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_5),
.B(n_321),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_5),
.B(n_362),
.Y(n_361)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_7),
.B(n_14),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_8),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_8),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_8),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_8),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_8),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_8),
.B(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_12),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_12),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_12),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_12),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_12),
.B(n_379),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_13),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_14),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_15),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_15),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_15),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_15),
.B(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_15),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_217),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_215),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_178),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_20),
.B(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.C(n_130),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_21),
.B(n_102),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_22),
.B(n_67),
.C(n_88),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_57),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_23),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_31),
.C(n_35),
.Y(n_101)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_26),
.Y(n_188)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_27),
.Y(n_157)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_30),
.A2(n_31),
.B1(n_235),
.B2(n_236),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_31),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_33),
.Y(n_338)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_34),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_35),
.A2(n_38),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_35),
.B(n_104),
.C(n_109),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_35),
.A2(n_38),
.B1(n_334),
.B2(n_339),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_35),
.B(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_37),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_39),
.B(n_57),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.C(n_50),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_41),
.B(n_51),
.Y(n_134)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_44),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_45),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_49),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_50),
.A2(n_51),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_55),
.Y(n_230)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_55),
.Y(n_295)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_56),
.Y(n_318)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_56),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_88),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_81),
.C(n_83),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_68),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.C(n_79),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_69),
.A2(n_70),
.B1(n_79),
.B2(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_69),
.A2(n_70),
.B1(n_117),
.B2(n_118),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_70),
.B(n_118),
.Y(n_266)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_73),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_73),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_74),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_78),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_101),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_100),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_90),
.A2(n_91),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_91),
.B(n_94),
.C(n_101),
.Y(n_203)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_98),
.Y(n_232)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_99),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_103),
.B(n_115),
.C(n_116),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_155),
.C(n_158),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_104),
.A2(n_112),
.B1(n_155),
.B2(n_258),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_106),
.Y(n_344)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_106),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_122),
.C(n_125),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_117),
.A2(n_118),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_129),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_130),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_161),
.C(n_175),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_131),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_153),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_133),
.B(n_154),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_135),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.C(n_149),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_136),
.A2(n_137),
.B1(n_149),
.B2(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_142),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_155),
.Y(n_258)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_175),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.C(n_171),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_162),
.B(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_162),
.A2(n_164),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_214),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_201),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_192),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_198),
.B2(n_200),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_229),
.C(n_231),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_198),
.A2(n_200),
.B1(n_231),
.B2(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_248),
.B(n_410),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_246),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_219),
.B(n_246),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_222),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_239),
.C(n_244),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_233),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_226),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_228),
.A2(n_233),
.B1(n_234),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_229),
.B(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_244),
.Y(n_254)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_306),
.B(n_406),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_277),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_251),
.A2(n_408),
.B(n_409),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_275),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_252),
.B(n_275),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.C(n_273),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_264),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_261),
.B(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_265),
.A2(n_266),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_304),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_278),
.B(n_304),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_301),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_279),
.B(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_281),
.B(n_301),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.C(n_299),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_282),
.B(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_285),
.A2(n_299),
.B1(n_300),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_285),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.C(n_296),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_286),
.A2(n_287),
.B1(n_296),
.B2(n_297),
.Y(n_385)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_291),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_401),
.B(n_405),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_387),
.B(n_400),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_374),
.B(n_386),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_350),
.B(n_373),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_340),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_340),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_325),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_326),
.C(n_333),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_319),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_313),
.B(n_320),
.C(n_322),
.Y(n_383)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_330),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_328),
.Y(n_362)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.C(n_345),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_345),
.B1(n_346),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_342),
.Y(n_371)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_367),
.B(n_372),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_360),
.B(n_366),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_359),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_359),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_357),
.Y(n_368)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_369),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_376),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_382),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_383),
.C(n_384),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_377),
.Y(n_411)
);

FAx1_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.CI(n_381),
.CON(n_377),
.SN(n_377)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_380),
.C(n_381),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_399),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_399),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_396),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_393),
.C(n_396),
.Y(n_402)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_403),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);


endmodule