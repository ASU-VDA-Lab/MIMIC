module fake_jpeg_19219_n_209 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_39),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_25),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_50),
.Y(n_56)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_53),
.B1(n_35),
.B2(n_49),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_57),
.B1(n_16),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_58),
.B(n_63),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_22),
.B(n_21),
.Y(n_61)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_65),
.B1(n_79),
.B2(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_16),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_26),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_30),
.B(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_30),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_23),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_92),
.C(n_108),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_102),
.B1(n_106),
.B2(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_111),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_15),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_71),
.Y(n_118)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_34),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_2),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_15),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_17),
.B1(n_15),
.B2(n_34),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_110),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_24),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_33),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_82),
.B1(n_59),
.B2(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_129),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_88),
.C(n_92),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_81),
.B1(n_74),
.B2(n_85),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_126),
.B1(n_94),
.B2(n_110),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_66),
.A3(n_81),
.B1(n_85),
.B2(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_130),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_60),
.C(n_59),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_127),
.C(n_114),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_106),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_4),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_146),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_109),
.B1(n_104),
.B2(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_143),
.B1(n_120),
.B2(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_101),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_99),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_130),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_102),
.C(n_103),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_105),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_123),
.B1(n_121),
.B2(n_113),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_122),
.B(n_134),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_136),
.B(n_149),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_149),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_134),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_139),
.B(n_145),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_120),
.B(n_89),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_154),
.B(n_137),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_148),
.C(n_151),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_141),
.C(n_153),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_139),
.C(n_140),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_162),
.B(n_158),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.C(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_168),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_136),
.Y(n_181)
);

OAI321xp33_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_164),
.B1(n_160),
.B2(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_157),
.B1(n_159),
.B2(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

FAx1_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_178),
.CI(n_170),
.CON(n_185),
.SN(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_168),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_173),
.B1(n_7),
.B2(n_9),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_177),
.B(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_6),
.C(n_7),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_174),
.C(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_9),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_185),
.B1(n_190),
.B2(n_197),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_202),
.B(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_10),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_10),
.Y(n_209)
);


endmodule