module fake_jpeg_15897_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_10),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_61),
.B1(n_57),
.B2(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_73),
.B1(n_48),
.B2(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_61),
.B1(n_54),
.B2(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_55),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_55),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_50),
.B(n_53),
.C(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_60),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_58),
.B1(n_48),
.B2(n_43),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_87),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_44),
.B1(n_48),
.B2(n_3),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_101),
.Y(n_111)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_89),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_96),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_1),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_97),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_24),
.B1(n_39),
.B2(n_38),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_70),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_7),
.Y(n_103)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_108),
.B1(n_95),
.B2(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_115),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_93),
.B1(n_108),
.B2(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_35),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_110),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_92),
.C(n_106),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_106),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_87),
.B1(n_109),
.B2(n_9),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_94),
.B1(n_107),
.B2(n_12),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_129),
.B1(n_124),
.B2(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_11),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_14),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_17),
.B(n_20),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_21),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_26),
.B(n_27),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_28),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_30),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_34),
.Y(n_141)
);


endmodule