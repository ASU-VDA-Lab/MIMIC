module real_jpeg_5634_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_0),
.A2(n_36),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_0),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_0),
.A2(n_256),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_0),
.A2(n_111),
.B1(n_256),
.B2(n_348),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_0),
.A2(n_88),
.B1(n_256),
.B2(n_441),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_1),
.A2(n_79),
.B1(n_177),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_1),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_287),
.C(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_1),
.B(n_75),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_1),
.B(n_159),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_1),
.B(n_124),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_1),
.B(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_2),
.A2(n_34),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_2),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_2),
.A2(n_112),
.B1(n_191),
.B2(n_283),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_2),
.A2(n_120),
.B1(n_160),
.B2(n_191),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_2),
.A2(n_191),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_3),
.Y(n_239)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_3),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_4),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_73),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_5),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_58),
.B1(n_90),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_90),
.B1(n_105),
.B2(n_181),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_90),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_6),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_7),
.A2(n_177),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_7),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_7),
.A2(n_307),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_7),
.A2(n_307),
.B1(n_396),
.B2(n_397),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_7),
.A2(n_33),
.B1(n_307),
.B2(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_8),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_35),
.B1(n_50),
.B2(n_53),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_53),
.B1(n_89),
.B2(n_200),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_9),
.A2(n_53),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_9),
.A2(n_53),
.B1(n_165),
.B2(n_294),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_10),
.Y(n_529)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_33),
.B1(n_57),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_12),
.A2(n_60),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_60),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_12),
.A2(n_60),
.B1(n_294),
.B2(n_315),
.Y(n_426)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_35),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_14),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_14),
.A2(n_186),
.B1(n_248),
.B2(n_252),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_14),
.A2(n_186),
.B1(n_234),
.B2(n_370),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_14),
.A2(n_186),
.B1(n_445),
.B2(n_448),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_15),
.Y(n_168)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_18),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_18),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_18),
.A2(n_98),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_18),
.A2(n_98),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_18),
.A2(n_98),
.B1(n_165),
.B2(n_169),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_524),
.B(n_526),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_147),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_145),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_141),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_23),
.B(n_141),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_131),
.C(n_138),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_24),
.A2(n_25),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_99),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_26),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_54),
.B1(n_56),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_27),
.A2(n_54),
.B1(n_132),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_27),
.A2(n_49),
.B1(n_54),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_27),
.A2(n_255),
.B(n_259),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_27),
.A2(n_54),
.B1(n_255),
.B2(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_28),
.B(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_28),
.A2(n_433),
.B(n_437),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_40),
.B1(n_43),
.B2(n_47),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_34),
.Y(n_143)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_41),
.B(n_354),
.Y(n_417)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_44),
.Y(n_364)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_45),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_46),
.Y(n_355)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_48),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_54),
.B(n_280),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_54),
.A2(n_189),
.B(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_55),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_55),
.B(n_190),
.Y(n_259)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_59),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_61),
.A2(n_99),
.B1(n_100),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_62),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_62),
.A2(n_87),
.B1(n_91),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_62),
.A2(n_91),
.B1(n_199),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_62),
.A2(n_91),
.B1(n_395),
.B2(n_440),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_75),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_73),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_68),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_73),
.Y(n_397)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_75),
.A2(n_139),
.B1(n_198),
.B2(n_203),
.Y(n_197)
);

AOI22x1_ASAP7_75t_L g471 ( 
.A1(n_75),
.A2(n_139),
.B1(n_399),
.B2(n_472),
.Y(n_471)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_78),
.Y(n_378)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_81),
.Y(n_245)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_81),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_81),
.Y(n_381)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_84),
.Y(n_450)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_91),
.B(n_362),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_91),
.A2(n_395),
.B(n_398),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_94),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_94),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_95),
.Y(n_396)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_99),
.A2(n_100),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_99),
.B(n_210),
.C(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_123),
.B(n_125),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_101),
.A2(n_279),
.B(n_281),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_101),
.A2(n_123),
.B1(n_304),
.B2(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_101),
.A2(n_281),
.B(n_347),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_101),
.A2(n_123),
.B1(n_444),
.B2(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_102),
.A2(n_124),
.B1(n_172),
.B2(n_180),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_102),
.A2(n_124),
.B1(n_180),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_102),
.A2(n_124),
.B1(n_172),
.B2(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_102),
.B(n_282),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_105),
.B(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_108),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_113),
.A2(n_304),
.B(n_308),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_120),
.B2(n_122),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_119),
.Y(n_370)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_123),
.A2(n_308),
.B(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_124),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_131),
.B(n_138),
.Y(n_521)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_136),
.Y(n_413)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_137),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_139),
.A2(n_352),
.B(n_361),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_139),
.B(n_399),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_139),
.A2(n_361),
.B(n_488),
.Y(n_487)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_144),
.B(n_280),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_518),
.B(n_523),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_271),
.B(n_515),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_260),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_217),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_151),
.B(n_217),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_151),
.Y(n_531)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_194),
.CI(n_208),
.CON(n_151),
.SN(n_151)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_152),
.B(n_194),
.C(n_208),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_183),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_171),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_154),
.A2(n_183),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_154),
.A2(n_171),
.B1(n_222),
.B2(n_459),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_163),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_155),
.A2(n_164),
.B1(n_229),
.B2(n_237),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_155),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_155),
.A2(n_280),
.B(n_297),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_155),
.A2(n_421),
.B1(n_422),
.B2(n_425),
.Y(n_420)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_156),
.B(n_300),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_156),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_156),
.A2(n_158),
.B1(n_369),
.B2(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_156),
.A2(n_298),
.B1(n_426),
.B2(n_465),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_168),
.Y(n_325)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_171),
.Y(n_459)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI32xp33_ASAP7_75t_L g371 ( 
.A1(n_174),
.A2(n_357),
.A3(n_372),
.B1(n_376),
.B2(n_379),
.Y(n_371)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g412 ( 
.A1(n_200),
.A2(n_413),
.A3(n_414),
.B1(n_417),
.B2(n_418),
.Y(n_412)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_216),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_210),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_209),
.B(n_262),
.C(n_266),
.Y(n_522)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.C(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_223),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_226),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_246),
.C(n_254),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_227),
.B(n_457),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_240),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_228),
.B(n_240),
.Y(n_482)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_229),
.Y(n_465)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_237),
.A2(n_320),
.B(n_326),
.Y(n_319)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_241),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_245),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_246),
.B(n_254),
.Y(n_457)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_247),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_253),
.Y(n_375)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_259),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_260),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_270),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_261),
.B(n_270),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI311xp33_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_453),
.A3(n_491),
.B1(n_509),
.C1(n_510),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_406),
.B(n_452),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_386),
.B(n_405),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_341),
.B(n_385),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_311),
.B(n_340),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_290),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_277),
.B(n_290),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_278),
.A2(n_284),
.B1(n_285),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_280),
.A2(n_353),
.B(n_356),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_SL g433 ( 
.A1(n_280),
.A2(n_418),
.B(n_434),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_301),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_302),
.C(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_299),
.A2(n_326),
.B(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_309),
.B2(n_310),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_329),
.B(n_339),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_318),
.B(n_328),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_327),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_327),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_337),
.Y(n_339)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_336),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_343),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_366),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_350),
.B2(n_351),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_350),
.C(n_366),
.Y(n_387)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_371),
.Y(n_392)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_387),
.B(n_388),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_393),
.B2(n_404),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_392),
.C(n_404),
.Y(n_407)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_400),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_401),
.C(n_402),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_407),
.B(n_408),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_430),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_409)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_419),
.B2(n_420),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_412),
.B(n_419),
.Y(n_486)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_427),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_428),
.C(n_430),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_438),
.B2(n_451),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_431),
.B(n_439),
.C(n_443),
.Y(n_500)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_443),
.Y(n_438)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_440),
.Y(n_488)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_476),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_SL g510 ( 
.A1(n_454),
.A2(n_476),
.B(n_511),
.C(n_514),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_473),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_455),
.B(n_473),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_460),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_458),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_466),
.C(n_471),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_464),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_466),
.A2(n_467),
.B1(n_471),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_471),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_489),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_489),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_482),
.C(n_483),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_486),
.C(n_487),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_484),
.A2(n_485),
.B1(n_487),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_487),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_504),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_493),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

NOR2x1_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_501),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_501),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_498),
.C(n_500),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_507),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_498),
.A2(n_499),
.B1(n_500),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_500),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_506),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_522),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_522),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx8_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);


endmodule