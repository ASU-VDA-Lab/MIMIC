module fake_jpeg_9541_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_41),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_48),
.B1(n_55),
.B2(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_40),
.B(n_31),
.C(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_41),
.B1(n_33),
.B2(n_19),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_63),
.B(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_22),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_33),
.C(n_28),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_16),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_43),
.B1(n_51),
.B2(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_23),
.B(n_39),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_96),
.B(n_23),
.Y(n_101)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_97),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_15),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_0),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_103),
.B(n_24),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_66),
.C(n_64),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_108),
.C(n_28),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_51),
.B1(n_92),
.B2(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_15),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_30),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_90),
.B1(n_81),
.B2(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_96),
.B1(n_94),
.B2(n_85),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_126),
.B(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_88),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_134),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_98),
.B1(n_94),
.B2(n_86),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_95),
.B1(n_93),
.B2(n_86),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_57),
.B(n_87),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_11),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_28),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_103),
.B(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_115),
.B(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_135),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_111),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_149),
.C(n_128),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_151),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_126),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_145),
.B(n_137),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_150),
.C(n_140),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_112),
.B1(n_116),
.B2(n_134),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_57),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_165),
.Y(n_174)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_57),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_170),
.C(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_140),
.C(n_145),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_166),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_144),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_177),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_157),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_174),
.C(n_160),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_185),
.Y(n_193)
);

OAI31xp33_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_154),
.A3(n_155),
.B(n_158),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_173),
.A3(n_156),
.B1(n_174),
.B2(n_12),
.C1(n_14),
.C2(n_8),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_192),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_182),
.B(n_180),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_12),
.B(n_2),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_188),
.B(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_1),
.C(n_2),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_194),
.A2(n_52),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_197),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_186),
.B(n_3),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_52),
.C(n_24),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_1),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_52),
.C2(n_202),
.Y(n_204)
);

NOR4xp25_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.C(n_6),
.D(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_6),
.Y(n_206)
);


endmodule