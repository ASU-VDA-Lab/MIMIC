module fake_jpeg_19962_n_67 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_25),
.B1(n_3),
.B2(n_5),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_45)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_15),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_28),
.C(n_9),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.C(n_43),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_8),
.C(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_52),
.B1(n_50),
.B2(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_64),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_17),
.C(n_20),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_22),
.Y(n_67)
);


endmodule