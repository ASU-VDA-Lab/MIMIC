module real_aes_8259_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_449;
wire n_417;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_0), .A2(n_208), .B(n_211), .C(n_292), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_1), .A2(n_241), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_2), .B(n_308), .Y(n_327) );
INVx1_ASAP7_75t_L g194 ( .A(n_3), .Y(n_194) );
AND2x6_ASAP7_75t_L g208 ( .A(n_3), .B(n_192), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_3), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g282 ( .A(n_4), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_5), .B(n_219), .Y(n_294) );
AOI22xp5_ASAP7_75t_SL g523 ( .A1(n_5), .A2(n_80), .B1(n_81), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_5), .Y(n_524) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_6), .A2(n_22), .B1(n_89), .B2(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g227 ( .A(n_7), .Y(n_227) );
INVx1_ASAP7_75t_L g152 ( .A(n_8), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_9), .A2(n_217), .B(n_304), .C(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_10), .B(n_308), .Y(n_307) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_11), .A2(n_24), .B1(n_89), .B2(n_90), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_12), .B(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_13), .A2(n_322), .B(n_337), .C(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_14), .B(n_219), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_15), .B(n_219), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_16), .Y(n_258) );
INVx1_ASAP7_75t_L g215 ( .A(n_17), .Y(n_215) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_18), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_19), .Y(n_290) );
INVx1_ASAP7_75t_L g247 ( .A(n_20), .Y(n_247) );
INVx2_ASAP7_75t_L g206 ( .A(n_21), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_23), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g185 ( .A1(n_24), .A2(n_43), .B1(n_55), .B2(n_186), .C(n_187), .Y(n_185) );
INVxp67_ASAP7_75t_L g188 ( .A(n_24), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_25), .A2(n_322), .B(n_323), .C(n_325), .Y(n_321) );
INVxp67_ASAP7_75t_L g248 ( .A(n_26), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_27), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g178 ( .A(n_27), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_28), .A2(n_211), .B(n_214), .C(n_222), .Y(n_210) );
CKINVDCx14_ASAP7_75t_R g320 ( .A(n_29), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_30), .A2(n_266), .B(n_280), .C(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g157 ( .A(n_31), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_32), .A2(n_80), .B1(n_81), .B2(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_32), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_33), .A2(n_174), .B1(n_175), .B2(n_179), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_33), .Y(n_174) );
INVx1_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_35), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_36), .Y(n_243) );
INVx1_ASAP7_75t_L g150 ( .A(n_37), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_38), .A2(n_39), .B1(n_84), .B2(n_100), .Y(n_83) );
AOI222xp33_ASAP7_75t_L g162 ( .A1(n_40), .A2(n_52), .B1(n_53), .B2(n_163), .C1(n_164), .C2(n_168), .Y(n_162) );
INVx1_ASAP7_75t_L g335 ( .A(n_41), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_42), .A2(n_173), .B1(n_180), .B2(n_181), .Y(n_172) );
INVx1_ASAP7_75t_L g180 ( .A(n_42), .Y(n_180) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_43), .A2(n_66), .B1(n_89), .B2(n_90), .Y(n_88) );
INVxp67_ASAP7_75t_L g189 ( .A(n_43), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_44), .A2(n_75), .B1(n_106), .B2(n_113), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g278 ( .A(n_45), .Y(n_278) );
INVx1_ASAP7_75t_L g192 ( .A(n_46), .Y(n_192) );
INVx1_ASAP7_75t_L g226 ( .A(n_47), .Y(n_226) );
INVx1_ASAP7_75t_L g119 ( .A(n_48), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_49), .Y(n_186) );
INVx1_ASAP7_75t_SL g324 ( .A(n_50), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_51), .B(n_308), .Y(n_340) );
INVx1_ASAP7_75t_L g261 ( .A(n_54), .Y(n_261) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_55), .A2(n_71), .B1(n_89), .B2(n_94), .Y(n_93) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_56), .A2(n_72), .B1(n_131), .B2(n_136), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_57), .A2(n_241), .B(n_277), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_58), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_59), .A2(n_241), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_60), .B(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_61), .A2(n_240), .B(n_242), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_62), .Y(n_209) );
INVx1_ASAP7_75t_L g302 ( .A(n_63), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_64), .A2(n_241), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g305 ( .A(n_65), .Y(n_305) );
INVx2_ASAP7_75t_L g224 ( .A(n_67), .Y(n_224) );
INVx1_ASAP7_75t_L g293 ( .A(n_68), .Y(n_293) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_69), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_70), .A2(n_211), .B(n_260), .C(n_268), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_73), .B(n_231), .Y(n_283) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_76), .A2(n_80), .B1(n_81), .B2(n_171), .Y(n_79) );
INVx2_ASAP7_75t_L g171 ( .A(n_76), .Y(n_171) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_182), .B1(n_195), .B2(n_519), .C(n_522), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_172), .Y(n_78) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND4xp75_ASAP7_75t_L g81 ( .A(n_82), .B(n_118), .C(n_140), .D(n_162), .Y(n_81) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_105), .Y(n_82) );
BUFx2_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x6_ASAP7_75t_L g156 ( .A(n_86), .B(n_128), .Y(n_156) );
AND2x4_ASAP7_75t_L g161 ( .A(n_86), .B(n_112), .Y(n_161) );
AND2x6_ASAP7_75t_L g163 ( .A(n_86), .B(n_139), .Y(n_163) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g104 ( .A(n_87), .B(n_93), .Y(n_104) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g110 ( .A(n_88), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_88), .B(n_93), .Y(n_117) );
AND2x2_ASAP7_75t_L g135 ( .A(n_88), .B(n_97), .Y(n_135) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g111 ( .A(n_93), .Y(n_111) );
INVx1_ASAP7_75t_L g167 ( .A(n_93), .Y(n_167) );
AND2x4_ASAP7_75t_L g103 ( .A(n_95), .B(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_95), .B(n_110), .Y(n_145) );
AND2x4_ASAP7_75t_L g148 ( .A(n_95), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g112 ( .A(n_96), .B(n_99), .Y(n_112) );
OR2x2_ASAP7_75t_L g129 ( .A(n_96), .B(n_99), .Y(n_129) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g139 ( .A(n_97), .B(n_99), .Y(n_139) );
AND2x2_ASAP7_75t_L g166 ( .A(n_98), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
INVx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx4_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2x1p5_ASAP7_75t_L g122 ( .A(n_104), .B(n_112), .Y(n_122) );
AND2x4_ASAP7_75t_L g127 ( .A(n_104), .B(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g138 ( .A(n_111), .Y(n_138) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx6_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OR2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx1_ASAP7_75t_L g134 ( .A(n_116), .Y(n_134) );
INVx1_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
OA211x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B(n_123), .C(n_130), .Y(n_118) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g165 ( .A(n_135), .B(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g169 ( .A(n_135), .B(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_151), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_146), .B2(n_150), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVxp67_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B1(n_157), .B2(n_158), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx11_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx6_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g170 ( .A(n_167), .Y(n_170) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_171), .B(n_249), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_173), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_175), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
AND3x1_ASAP7_75t_SL g184 ( .A(n_185), .B(n_190), .C(n_193), .Y(n_184) );
INVxp67_ASAP7_75t_L g528 ( .A(n_185), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_SL g529 ( .A(n_190), .Y(n_529) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_190), .A2(n_204), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g539 ( .A(n_190), .Y(n_539) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_191), .B(n_194), .Y(n_533) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_SL g538 ( .A(n_193), .B(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR4x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_409), .C(n_456), .D(n_496), .Y(n_196) );
NAND3xp33_ASAP7_75t_SL g197 ( .A(n_198), .B(n_355), .C(n_384), .Y(n_197) );
AOI211xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_271), .B(n_309), .C(n_348), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_199), .A2(n_368), .B(n_385), .C(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_233), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_201), .B(n_347), .Y(n_346) );
INVx3_ASAP7_75t_SL g351 ( .A(n_201), .Y(n_351) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_201), .Y(n_363) );
AND2x4_ASAP7_75t_L g367 ( .A(n_201), .B(n_316), .Y(n_367) );
AND2x2_ASAP7_75t_L g378 ( .A(n_201), .B(n_256), .Y(n_378) );
OR2x2_ASAP7_75t_L g402 ( .A(n_201), .B(n_312), .Y(n_402) );
AND2x2_ASAP7_75t_L g415 ( .A(n_201), .B(n_317), .Y(n_415) );
AND2x2_ASAP7_75t_L g455 ( .A(n_201), .B(n_441), .Y(n_455) );
AND2x2_ASAP7_75t_L g462 ( .A(n_201), .B(n_425), .Y(n_462) );
AND2x2_ASAP7_75t_L g492 ( .A(n_201), .B(n_234), .Y(n_492) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_228), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_209), .B(n_210), .C(n_223), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_203), .A2(n_258), .B(n_259), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_203), .A2(n_290), .B(n_291), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_204), .B(n_208), .Y(n_203) );
AND2x4_ASAP7_75t_L g241 ( .A(n_204), .B(n_208), .Y(n_241) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
INVx1_ASAP7_75t_L g221 ( .A(n_205), .Y(n_221) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g212 ( .A(n_206), .Y(n_212) );
INVx1_ASAP7_75t_L g339 ( .A(n_206), .Y(n_339) );
INVx1_ASAP7_75t_L g213 ( .A(n_207), .Y(n_213) );
INVx3_ASAP7_75t_L g217 ( .A(n_207), .Y(n_217) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_207), .Y(n_219) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_207), .Y(n_250) );
BUFx3_ASAP7_75t_L g222 ( .A(n_208), .Y(n_222) );
INVx4_ASAP7_75t_SL g251 ( .A(n_208), .Y(n_251) );
INVx5_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
AND2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
BUFx3_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_212), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_218), .C(n_220), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_216), .A2(n_247), .B1(n_248), .B2(n_249), .Y(n_246) );
INVx5_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_217), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
INVx4_ASAP7_75t_L g322 ( .A(n_219), .Y(n_322) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_221), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g254 ( .A(n_223), .Y(n_254) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_223), .A2(n_276), .B(n_283), .Y(n_275) );
INVx1_ASAP7_75t_L g288 ( .A(n_223), .Y(n_288) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_L g232 ( .A(n_224), .B(n_225), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_230), .A2(n_257), .B(n_269), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_230), .B(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g238 ( .A(n_232), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_233), .B(n_419), .Y(n_431) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_255), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_234), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g369 ( .A(n_234), .B(n_255), .Y(n_369) );
BUFx3_ASAP7_75t_L g377 ( .A(n_234), .Y(n_377) );
OR2x2_ASAP7_75t_L g398 ( .A(n_234), .B(n_274), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_234), .B(n_419), .Y(n_509) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_239), .B(n_252), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_236), .A2(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_240), .Y(n_521) );
BUFx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_243), .A2(n_244), .B(n_245), .C(n_251), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g277 ( .A1(n_244), .A2(n_251), .B(n_278), .C(n_279), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_SL g301 ( .A1(n_244), .A2(n_251), .B(n_302), .C(n_303), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_244), .A2(n_251), .B(n_320), .C(n_321), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_SL g334 ( .A1(n_244), .A2(n_251), .B(n_335), .C(n_336), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_249), .B(n_305), .Y(n_304) );
INVx4_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g263 ( .A(n_250), .Y(n_263) );
INVx1_ASAP7_75t_L g268 ( .A(n_251), .Y(n_268) );
INVx1_ASAP7_75t_L g314 ( .A(n_252), .Y(n_314) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_254), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g315 ( .A(n_255), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g362 ( .A(n_255), .Y(n_362) );
AND2x2_ASAP7_75t_L g425 ( .A(n_255), .B(n_317), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_255), .A2(n_428), .B1(n_430), .B2(n_432), .C(n_433), .Y(n_427) );
AND2x2_ASAP7_75t_L g441 ( .A(n_255), .B(n_312), .Y(n_441) );
AND2x2_ASAP7_75t_L g467 ( .A(n_255), .B(n_351), .Y(n_467) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g347 ( .A(n_256), .B(n_317), .Y(n_347) );
BUFx2_ASAP7_75t_L g481 ( .A(n_256), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_264), .C(n_265), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_L g292 ( .A1(n_262), .A2(n_265), .B(n_293), .C(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI32xp33_ASAP7_75t_L g447 ( .A1(n_272), .A2(n_408), .A3(n_422), .B1(n_448), .B2(n_449), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_284), .Y(n_272) );
AND2x2_ASAP7_75t_L g388 ( .A(n_273), .B(n_331), .Y(n_388) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g370 ( .A(n_274), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_274), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g442 ( .A(n_274), .B(n_331), .Y(n_442) );
AND2x2_ASAP7_75t_L g453 ( .A(n_274), .B(n_345), .Y(n_453) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g354 ( .A(n_275), .B(n_332), .Y(n_354) );
AND2x2_ASAP7_75t_L g358 ( .A(n_275), .B(n_332), .Y(n_358) );
AND2x2_ASAP7_75t_L g393 ( .A(n_275), .B(n_344), .Y(n_393) );
AND2x2_ASAP7_75t_L g400 ( .A(n_275), .B(n_297), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_275), .A2(n_351), .B(n_362), .C(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g459 ( .A(n_275), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_275), .B(n_286), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_284), .B(n_342), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_284), .B(n_358), .Y(n_448) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g353 ( .A(n_285), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_297), .Y(n_285) );
AND2x2_ASAP7_75t_L g345 ( .A(n_286), .B(n_298), .Y(n_345) );
OR2x2_ASAP7_75t_L g360 ( .A(n_286), .B(n_298), .Y(n_360) );
AND2x2_ASAP7_75t_L g383 ( .A(n_286), .B(n_344), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_286), .Y(n_387) );
AND2x2_ASAP7_75t_L g406 ( .A(n_286), .B(n_343), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_286), .A2(n_371), .B1(n_417), .B2(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_286), .B(n_459), .Y(n_483) );
AND2x2_ASAP7_75t_L g498 ( .A(n_286), .B(n_358), .Y(n_498) );
INVx4_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g329 ( .A(n_287), .Y(n_329) );
AND2x2_ASAP7_75t_L g372 ( .A(n_287), .B(n_298), .Y(n_372) );
AND2x2_ASAP7_75t_L g374 ( .A(n_287), .B(n_331), .Y(n_374) );
AND3x2_ASAP7_75t_L g436 ( .A(n_287), .B(n_400), .C(n_437), .Y(n_436) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_295), .Y(n_287) );
OAI322xp33_ASAP7_75t_L g522 ( .A1(n_290), .A2(n_523), .A3(n_525), .B1(n_529), .B2(n_530), .C1(n_534), .C2(n_536), .Y(n_522) );
AND2x2_ASAP7_75t_L g471 ( .A(n_297), .B(n_343), .Y(n_471) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g331 ( .A(n_298), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_298), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_298), .B(n_342), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_298), .B(n_383), .C(n_459), .Y(n_511) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_307), .Y(n_298) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_299), .A2(n_318), .B(n_327), .Y(n_317) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_299), .A2(n_333), .B(n_340), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_328), .B1(n_341), .B2(n_346), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_312), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g423 ( .A(n_312), .Y(n_423) );
OAI31xp33_ASAP7_75t_L g439 ( .A1(n_315), .A2(n_440), .A3(n_441), .B(n_442), .Y(n_439) );
AND2x2_ASAP7_75t_L g464 ( .A(n_315), .B(n_351), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_315), .B(n_377), .Y(n_510) );
AND2x2_ASAP7_75t_L g419 ( .A(n_316), .B(n_351), .Y(n_419) );
AND2x2_ASAP7_75t_L g480 ( .A(n_316), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g408 ( .A(n_317), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_322), .B(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_329), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_330), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AOI221x1_ASAP7_75t_SL g396 ( .A1(n_331), .A2(n_397), .B1(n_399), .B2(n_401), .C(n_403), .Y(n_396) );
INVx2_ASAP7_75t_L g344 ( .A(n_332), .Y(n_344) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_332), .Y(n_438) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g426 ( .A(n_341), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_342), .B(n_359), .Y(n_451) );
INVx1_ASAP7_75t_SL g514 ( .A(n_342), .Y(n_514) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g432 ( .A(n_345), .B(n_358), .Y(n_432) );
INVx1_ASAP7_75t_L g500 ( .A(n_346), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_346), .B(n_429), .Y(n_513) );
INVx2_ASAP7_75t_SL g352 ( .A(n_347), .Y(n_352) );
AND2x2_ASAP7_75t_L g395 ( .A(n_347), .B(n_351), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_347), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_347), .B(n_422), .Y(n_449) );
AOI21xp33_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_352), .B(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_350), .B(n_422), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_350), .B(n_377), .Y(n_518) );
OR2x2_ASAP7_75t_L g390 ( .A(n_351), .B(n_369), .Y(n_390) );
AND2x2_ASAP7_75t_L g489 ( .A(n_351), .B(n_480), .Y(n_489) );
OAI22xp5_ASAP7_75t_SL g364 ( .A1(n_352), .A2(n_365), .B1(n_370), .B2(n_373), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_352), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g412 ( .A(n_354), .B(n_360), .Y(n_412) );
INVx1_ASAP7_75t_L g476 ( .A(n_354), .Y(n_476) );
AOI311xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .A3(n_363), .B(n_364), .C(n_375), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_359), .A2(n_491), .B1(n_503), .B2(n_506), .C(n_508), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_359), .B(n_514), .Y(n_516) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g413 ( .A(n_361), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g403 ( .A1(n_362), .A2(n_404), .B(n_405), .C(n_407), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_366), .A2(n_368), .B(n_473), .C(n_474), .Y(n_472) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_367), .B(n_441), .Y(n_507) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_370), .A2(n_390), .B1(n_391), .B2(n_394), .C(n_396), .Y(n_389) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g392 ( .A(n_372), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g475 ( .A(n_372), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_379), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_376), .A2(n_434), .B(n_435), .C(n_439), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_377), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_377), .B(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g399 ( .A(n_383), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_387), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g501 ( .A(n_390), .Y(n_501) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_393), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g428 ( .A(n_393), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g505 ( .A(n_393), .Y(n_505) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g446 ( .A(n_395), .B(n_422), .Y(n_446) );
INVx1_ASAP7_75t_SL g440 ( .A(n_402), .Y(n_440) );
INVx1_ASAP7_75t_L g417 ( .A(n_408), .Y(n_417) );
NAND3xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_427), .C(n_443), .Y(n_409) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .A3(n_414), .B1(n_416), .B2(n_420), .C1(n_424), .C2(n_426), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_411), .A2(n_464), .B(n_465), .C(n_472), .Y(n_463) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_414), .A2(n_435), .B1(n_466), .B2(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g424 ( .A(n_422), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g461 ( .A(n_422), .B(n_462), .Y(n_461) );
AOI32xp33_ASAP7_75t_L g512 ( .A1(n_422), .A2(n_513), .A3(n_514), .B1(n_515), .B2(n_517), .Y(n_512) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g434 ( .A(n_425), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_425), .A2(n_478), .B1(n_482), .B2(n_484), .C(n_487), .Y(n_477) );
AND2x2_ASAP7_75t_L g491 ( .A(n_425), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g494 ( .A(n_429), .B(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g504 ( .A(n_429), .B(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g495 ( .A(n_438), .B(n_459), .Y(n_495) );
AOI211xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B(n_447), .C(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_460), .B(n_463), .C(n_477), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_471), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_483), .Y(n_486) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_493), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI211xp5_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_499), .B(n_502), .C(n_512), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
endmodule