module fake_jpeg_13248_n_185 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_16),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_27),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_92),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_94),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_62),
.C(n_68),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_0),
.B(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_65),
.B1(n_86),
.B2(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_111),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_65),
.B1(n_86),
.B2(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_70),
.B1(n_59),
.B2(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_58),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_57),
.B1(n_81),
.B2(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_81),
.B1(n_80),
.B2(n_83),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_14),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_113)
);

AO22x2_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_75),
.B1(n_79),
.B2(n_76),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_75),
.C(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_125),
.Y(n_142)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_131),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_78),
.B1(n_73),
.B2(n_72),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_141)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_66),
.B1(n_64),
.B2(n_61),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_15),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_71),
.B1(n_5),
.B2(n_6),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_71),
.B1(n_26),
.B2(n_28),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_22),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_8),
.C(n_9),
.Y(n_135)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_6),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_138),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_29),
.C(n_53),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_24),
.C(n_52),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_140),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_146),
.B(n_123),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_33),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_54),
.B1(n_43),
.B2(n_45),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_14),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_15),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_130),
.B(n_17),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_32),
.B(n_35),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_39),
.B(n_47),
.C(n_48),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_158),
.C(n_153),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.C(n_142),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_156),
.B1(n_150),
.B2(n_152),
.C(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_174),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_175),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_169),
.B(n_168),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_166),
.C(n_159),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_134),
.C(n_171),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_158),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_140),
.Y(n_185)
);


endmodule