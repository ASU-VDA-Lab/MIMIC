module fake_netlist_1_9177_n_739 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_739);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_739;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_55), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_61), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_74), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_78), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_52), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_27), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_43), .Y(n_87) );
INVx3_ASAP7_75t_L g88 ( .A(n_9), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_7), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_16), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_51), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_11), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_9), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_76), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_53), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_80), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_50), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_41), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_31), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_73), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_26), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_30), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_58), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_32), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_79), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_35), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_70), .Y(n_125) );
INVxp33_ASAP7_75t_L g126 ( .A(n_14), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_13), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_98), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_116), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_81), .B(n_28), .Y(n_135) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_88), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_82), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_89), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_114), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_122), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_110), .Y(n_145) );
NOR2xp33_ASAP7_75t_R g146 ( .A(n_117), .B(n_29), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_81), .B(n_0), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_89), .B(n_1), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
NAND2xp33_ASAP7_75t_R g150 ( .A(n_125), .B(n_33), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_95), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
NOR2xp33_ASAP7_75t_SL g153 ( .A(n_124), .B(n_34), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_92), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_83), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_86), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_85), .B(n_2), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_93), .B(n_3), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_94), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_96), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_96), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_99), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_97), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_99), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_100), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_97), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_100), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_101), .Y(n_172) );
INVxp67_ASAP7_75t_L g173 ( .A(n_106), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_106), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
AO22x2_ASAP7_75t_L g180 ( .A1(n_148), .A2(n_130), .B1(n_129), .B2(n_101), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_155), .B(n_130), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_134), .B(n_136), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_148), .A2(n_111), .B1(n_128), .B2(n_113), .Y(n_196) );
OAI221xp5_ASAP7_75t_L g197 ( .A1(n_173), .A2(n_111), .B1(n_128), .B2(n_113), .C(n_115), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_138), .B(n_129), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_161), .B(n_115), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_138), .B(n_123), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_142), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_149), .B(n_90), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
CKINVDCx8_ASAP7_75t_R g211 ( .A(n_132), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_140), .B(n_123), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_166), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_160), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_166), .B(n_121), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_162), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_168), .B(n_121), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_168), .B(n_120), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_172), .B(n_107), .Y(n_226) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_147), .B(n_159), .C(n_139), .Y(n_227) );
OR2x6_ASAP7_75t_L g228 ( .A(n_164), .B(n_120), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_172), .B(n_119), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_167), .B(n_119), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_164), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_156), .B(n_118), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_169), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_140), .B(n_118), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_169), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_170), .Y(n_236) );
INVx4_ASAP7_75t_L g237 ( .A(n_157), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_154), .Y(n_238) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_141), .A2(n_104), .B1(n_91), .B2(n_103), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
AND2x6_ASAP7_75t_L g241 ( .A(n_150), .B(n_112), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_163), .B(n_112), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
INVx4_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_182), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
AND2x6_ASAP7_75t_SL g247 ( .A(n_202), .B(n_151), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_189), .B(n_146), .Y(n_248) );
NAND2xp33_ASAP7_75t_SL g249 ( .A(n_237), .B(n_174), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_211), .B(n_174), .Y(n_250) );
NOR2xp33_ASAP7_75t_R g251 ( .A(n_211), .B(n_165), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
INVxp67_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_200), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_189), .B(n_165), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_212), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_176), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
NOR2xp33_ASAP7_75t_R g262 ( .A(n_212), .B(n_163), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_176), .Y(n_263) );
INVx3_ASAP7_75t_SL g264 ( .A(n_237), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
NOR2xp33_ASAP7_75t_R g266 ( .A(n_176), .B(n_151), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_181), .B(n_3), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
INVx6_ASAP7_75t_L g269 ( .A(n_216), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_184), .B(n_109), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_224), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_235), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g275 ( .A(n_197), .B(n_4), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
NOR2xp33_ASAP7_75t_R g277 ( .A(n_181), .B(n_5), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
INVx5_ASAP7_75t_L g279 ( .A(n_228), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_181), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_227), .A2(n_105), .B1(n_87), .B2(n_107), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_180), .A2(n_109), .B1(n_108), .B2(n_102), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_189), .B(n_108), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_215), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_189), .B(n_102), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_209), .B(n_5), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_200), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_215), .B(n_6), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_183), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_196), .A2(n_6), .B1(n_8), .B2(n_10), .C(n_11), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_180), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_239), .B(n_8), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_180), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_188), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_217), .B(n_12), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_200), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_184), .B(n_39), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_221), .B(n_12), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_217), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_242), .B(n_13), .Y(n_307) );
NOR3xp33_ASAP7_75t_SL g308 ( .A(n_205), .B(n_14), .C(n_15), .Y(n_308) );
NOR3xp33_ASAP7_75t_SL g309 ( .A(n_214), .B(n_15), .C(n_16), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_232), .B(n_45), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_198), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_188), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_221), .B(n_17), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_221), .B(n_18), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_304), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_279), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_245), .B(n_239), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_279), .B(n_223), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
BUFx5_ASAP7_75t_L g323 ( .A(n_259), .Y(n_323) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
INVx3_ASAP7_75t_SL g326 ( .A(n_264), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_255), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
BUFx10_ASAP7_75t_L g329 ( .A(n_314), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_256), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_314), .A2(n_221), .B1(n_223), .B2(n_226), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_223), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_271), .A2(n_184), .B(n_187), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_261), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_265), .B(n_223), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_270), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_272), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_244), .B(n_226), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_297), .A2(n_215), .B1(n_180), .B2(n_198), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_262), .Y(n_341) );
CKINVDCx6p67_ASAP7_75t_R g342 ( .A(n_264), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_255), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_253), .B(n_226), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_250), .Y(n_345) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
BUFx10_ASAP7_75t_L g347 ( .A(n_278), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_271), .A2(n_184), .B(n_194), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_273), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_248), .B(n_226), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_286), .A2(n_194), .B(n_187), .Y(n_351) );
OR2x6_ASAP7_75t_L g352 ( .A(n_281), .B(n_204), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_291), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_299), .A2(n_234), .B1(n_225), .B2(n_229), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_255), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_258), .B(n_204), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_283), .B(n_236), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_287), .B(n_236), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_292), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_284), .B(n_204), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_278), .B(n_204), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_276), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_280), .B(n_299), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_301), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_290), .B(n_241), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_262), .B(n_185), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_280), .B(n_208), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_269), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_285), .A2(n_249), .B1(n_301), .B2(n_275), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_307), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_324), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_315), .B(n_198), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_319), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_326), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_335), .B(n_298), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_331), .B(n_294), .Y(n_377) );
INVx6_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_365), .A2(n_303), .B(n_305), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_324), .A2(n_250), .B1(n_251), .B2(n_266), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_332), .A2(n_296), .B1(n_311), .B2(n_208), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_311), .B1(n_198), .B2(n_208), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_369), .A2(n_294), .B1(n_313), .B2(n_208), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_350), .B(n_201), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_326), .B(n_230), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_363), .B(n_246), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_319), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_322), .Y(n_388) );
BUFx10_ASAP7_75t_L g389 ( .A(n_338), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_246), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_337), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_346), .A2(n_251), .B1(n_266), .B2(n_306), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_339), .A2(n_233), .A3(n_219), .B(n_220), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_346), .A2(n_277), .B1(n_267), .B2(n_241), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_303), .B(n_267), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_322), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_329), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_322), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_337), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_338), .B(n_289), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_320), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_322), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_360), .A2(n_309), .B1(n_308), .B2(n_241), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_382), .A2(n_359), .B1(n_366), .B2(n_317), .C(n_336), .Y(n_405) );
INVx6_ASAP7_75t_L g406 ( .A(n_389), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_382), .A2(n_356), .B1(n_352), .B2(n_338), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_391), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_371), .B(n_321), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_377), .A2(n_341), .B1(n_345), .B2(n_329), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_398), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_391), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_400), .B(n_330), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_404), .B(n_354), .C(n_310), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_377), .A2(n_356), .B1(n_345), .B2(n_361), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_403), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_377), .A2(n_329), .B1(n_356), .B2(n_277), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_371), .B(n_334), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_392), .A2(n_318), .B(n_361), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g423 ( .A1(n_392), .A2(n_352), .B1(n_247), .B2(n_318), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_404), .B(n_310), .C(n_353), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_402), .B(n_349), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_383), .A2(n_370), .B(n_355), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_394), .A2(n_352), .B1(n_357), .B2(n_358), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_318), .B(n_368), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_385), .A2(n_238), .B1(n_325), .B2(n_340), .C(n_289), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_388), .A2(n_370), .B(n_355), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_408), .B(n_393), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g436 ( .A1(n_423), .A2(n_381), .B1(n_380), .B2(n_375), .C1(n_372), .C2(n_384), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_423), .A2(n_342), .B1(n_375), .B2(n_381), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_405), .A2(n_376), .B1(n_384), .B2(n_373), .C(n_401), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_342), .B1(n_376), .B2(n_398), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_431), .B(n_398), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_409), .A2(n_401), .B1(n_201), .B2(n_203), .C(n_361), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_412), .B(n_374), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_422), .A2(n_394), .B(n_397), .C(n_398), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_421), .B(n_401), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_429), .A2(n_378), .B1(n_386), .B2(n_390), .Y(n_450) );
NOR2xp33_ASAP7_75t_R g451 ( .A(n_406), .B(n_378), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_416), .A2(n_401), .B1(n_390), .B2(n_386), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_426), .B(n_393), .Y(n_454) );
OR2x6_ASAP7_75t_L g455 ( .A(n_406), .B(n_378), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_411), .B(n_378), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
OAI33xp33_ASAP7_75t_L g459 ( .A1(n_414), .A2(n_190), .A3(n_191), .B1(n_192), .B2(n_195), .B3(n_193), .Y(n_459) );
OAI321xp33_ASAP7_75t_L g460 ( .A1(n_415), .A2(n_397), .A3(n_240), .B1(n_386), .B2(n_390), .C(n_368), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_430), .A2(n_401), .B1(n_203), .B2(n_397), .C(n_233), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_410), .A2(n_378), .B1(n_374), .B2(n_387), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_411), .B(n_374), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_411), .B(n_389), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_427), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_428), .B(n_393), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_433), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_428), .B(n_393), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_432), .B(n_389), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_454), .B(n_417), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_442), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_454), .B(n_427), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_457), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_468), .A2(n_427), .B(n_415), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_468), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_437), .B(n_389), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_436), .B(n_425), .C(n_420), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_469), .B(n_427), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_450), .A2(n_425), .B1(n_387), .B2(n_325), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_449), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_458), .A2(n_213), .B1(n_219), .B2(n_220), .C(n_231), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_434), .B(n_393), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g486 ( .A1(n_448), .A2(n_206), .A3(n_191), .B1(n_192), .B2(n_193), .B3(n_195), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_462), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_469), .B(n_393), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_462), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_438), .A2(n_241), .B1(n_387), .B2(n_395), .Y(n_490) );
OAI33xp33_ASAP7_75t_L g491 ( .A1(n_456), .A2(n_206), .A3(n_190), .B1(n_175), .B2(n_199), .B3(n_177), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_393), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_435), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_453), .B(n_417), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_453), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_467), .B(n_433), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_467), .B(n_433), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_445), .B(n_433), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_466), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_445), .B(n_418), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_447), .B(n_418), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_451), .Y(n_506) );
NAND2x1_ASAP7_75t_SL g507 ( .A(n_464), .B(n_388), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_464), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_464), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_457), .B(n_418), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_446), .B(n_175), .C(n_177), .Y(n_511) );
AOI21xp33_ASAP7_75t_SL g512 ( .A1(n_463), .A2(n_20), .B(n_22), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_418), .Y(n_513) );
AO221x2_ASAP7_75t_L g514 ( .A1(n_440), .A2(n_388), .B1(n_399), .B2(n_396), .C(n_395), .Y(n_514) );
OAI21xp5_ASAP7_75t_SL g515 ( .A1(n_439), .A2(n_340), .B(n_316), .Y(n_515) );
NAND4xp25_ASAP7_75t_SL g516 ( .A(n_444), .B(n_240), .C(n_231), .D(n_213), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_470), .A2(n_241), .B1(n_395), .B2(n_379), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_457), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_435), .B(n_419), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_443), .B(n_419), .Y(n_521) );
AOI21x1_ASAP7_75t_L g522 ( .A1(n_455), .A2(n_399), .B(n_396), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_455), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_455), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_478), .B(n_452), .C(n_461), .D(n_465), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_473), .B(n_419), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_495), .B(n_455), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_495), .B(n_419), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_472), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_475), .A2(n_459), .B(n_418), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_419), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_471), .B(n_451), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_487), .B(n_241), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_489), .B(n_396), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_471), .B(n_395), .Y(n_535) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_506), .B(n_328), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_471), .B(n_399), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_493), .B(n_241), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_471), .B(n_379), .Y(n_539) );
NAND2xp33_ASAP7_75t_R g540 ( .A(n_506), .B(n_460), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_498), .B(n_403), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_481), .B(n_379), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_494), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g546 ( .A(n_523), .B(n_474), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_494), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_504), .B(n_379), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_482), .Y(n_549) );
OR2x6_ASAP7_75t_L g550 ( .A(n_474), .B(n_403), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_520), .B(n_500), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_482), .Y(n_552) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_523), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_520), .B(n_347), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_476), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_485), .B(n_316), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_500), .B(n_347), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_508), .B(n_328), .Y(n_558) );
NOR2xp33_ASAP7_75t_R g559 ( .A(n_516), .B(n_316), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_485), .B(n_367), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_512), .B(n_24), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_498), .B(n_403), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_476), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_508), .B(n_36), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_509), .B(n_403), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_514), .A2(n_362), .B(n_343), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
INVx4_ASAP7_75t_L g568 ( .A(n_523), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_499), .B(n_199), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_488), .B(n_207), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_507), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_512), .B(n_179), .C(n_186), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_488), .B(n_367), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_477), .B(n_37), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_501), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_496), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_479), .B(n_367), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_484), .B(n_207), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_496), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_484), .B(n_210), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_511), .B(n_210), .C(n_186), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_503), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_576), .Y(n_587) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_525), .A2(n_515), .B(n_509), .C(n_518), .Y(n_588) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_574), .B(n_561), .C(n_577), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_572), .B(n_479), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_578), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_566), .A2(n_514), .B(n_491), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_529), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_542), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_543), .Y(n_595) );
OAI22xp33_ASAP7_75t_SL g596 ( .A1(n_545), .A2(n_474), .B1(n_518), .B2(n_524), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_577), .A2(n_490), .B(n_507), .C(n_517), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_540), .A2(n_561), .B1(n_546), .B2(n_568), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_540), .A2(n_546), .B1(n_568), .B2(n_553), .C(n_536), .Y(n_599) );
AOI32xp33_ASAP7_75t_L g600 ( .A1(n_547), .A2(n_480), .A3(n_524), .B1(n_510), .B2(n_513), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_566), .A2(n_514), .B(n_486), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_532), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_549), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_586), .B(n_492), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_530), .A2(n_514), .B(n_513), .Y(n_605) );
OA211x2_ASAP7_75t_L g606 ( .A1(n_568), .A2(n_522), .B(n_483), .C(n_521), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_563), .A2(n_505), .B(n_492), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_527), .B(n_503), .C(n_502), .D(n_510), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_563), .A2(n_505), .B1(n_502), .B2(n_519), .C(n_522), .Y(n_609) );
OAI31xp33_ASAP7_75t_L g610 ( .A1(n_557), .A2(n_519), .A3(n_521), .B(n_179), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_552), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_570), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_555), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_551), .B(n_521), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_579), .B(n_38), .Y(n_615) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_573), .A2(n_42), .B(n_44), .Y(n_616) );
OAI21xp33_ASAP7_75t_SL g617 ( .A1(n_573), .A2(n_46), .B(n_49), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_582), .B(n_54), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_539), .A2(n_323), .B1(n_269), .B2(n_268), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_571), .B(n_56), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_567), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_555), .B(n_60), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_571), .B(n_62), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_583), .B(n_63), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_530), .A2(n_362), .B(n_343), .Y(n_627) );
NOR2xp67_ASAP7_75t_SL g628 ( .A(n_585), .B(n_362), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_541), .B(n_64), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_548), .B(n_71), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_550), .A2(n_269), .B1(n_362), .B2(n_343), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_581), .A2(n_75), .B(n_77), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_575), .B(n_323), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_562), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_580), .B(n_323), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_556), .A2(n_351), .B(n_348), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_526), .B(n_343), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_526), .B(n_323), .Y(n_639) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_528), .A2(n_187), .A3(n_194), .B1(n_282), .B2(n_263), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_613), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_599), .A2(n_550), .B(n_544), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_641), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_589), .A2(n_531), .B1(n_539), .B2(n_535), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_614), .B(n_531), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_599), .B(n_533), .C(n_560), .Y(n_647) );
NAND2xp33_ASAP7_75t_R g648 ( .A(n_605), .B(n_559), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_590), .B(n_635), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_602), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_619), .B(n_537), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_622), .Y(n_652) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_596), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_633), .B(n_558), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_587), .Y(n_655) );
NAND2xp33_ASAP7_75t_L g656 ( .A(n_598), .B(n_559), .Y(n_656) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_600), .A2(n_550), .B1(n_538), .B2(n_564), .C(n_554), .Y(n_657) );
NOR3xp33_ASAP7_75t_SL g658 ( .A(n_597), .B(n_333), .C(n_565), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_608), .A2(n_565), .B(n_323), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_591), .Y(n_660) );
NAND2xp33_ASAP7_75t_L g661 ( .A(n_607), .B(n_565), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_588), .A2(n_609), .B(n_617), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_609), .B(n_323), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_604), .B(n_327), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_593), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_629), .Y(n_666) );
NOR3xp33_ASAP7_75t_SL g667 ( .A(n_616), .B(n_200), .C(n_327), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_624), .B(n_327), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_594), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_595), .B(n_243), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_603), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_611), .Y(n_672) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_610), .B(n_327), .C(n_243), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_623), .B(n_312), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_612), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_639), .B(n_312), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_638), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_630), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_605), .B(n_295), .Y(n_679) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_656), .B(n_601), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_659), .B(n_601), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_652), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_656), .A2(n_606), .B1(n_634), .B2(n_636), .Y(n_683) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_642), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_669), .B(n_621), .Y(n_685) );
NAND2x1_ASAP7_75t_L g686 ( .A(n_642), .B(n_627), .Y(n_686) );
XOR2xp5_ASAP7_75t_L g687 ( .A(n_645), .B(n_625), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_649), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_650), .A2(n_592), .B1(n_620), .B2(n_615), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_649), .B(n_592), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_644), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_672), .B(n_627), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_646), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_677), .B(n_618), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_648), .A2(n_626), .B1(n_632), .B2(n_631), .Y(n_695) );
OAI332xp33_ASAP7_75t_L g696 ( .A1(n_653), .A2(n_637), .A3(n_628), .B1(n_640), .B2(n_274), .B3(n_260), .C1(n_300), .C2(n_295), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_662), .A2(n_300), .B(n_260), .C(n_274), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_651), .B(n_259), .Y(n_698) );
OAI21xp5_ASAP7_75t_SL g699 ( .A1(n_643), .A2(n_276), .B(n_288), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_677), .B(n_276), .Y(n_700) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_654), .B(n_263), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_655), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_678), .B(n_282), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_703), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_691), .B(n_665), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_690), .B(n_666), .Y(n_706) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_680), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
NAND2xp33_ASAP7_75t_R g709 ( .A(n_692), .B(n_667), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_697), .A2(n_648), .B1(n_658), .B2(n_661), .C(n_657), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_688), .B(n_671), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_697), .B(n_679), .C(n_661), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_683), .A2(n_663), .B1(n_647), .B2(n_678), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_693), .A2(n_673), .B1(n_663), .B2(n_642), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_687), .A2(n_675), .B1(n_660), .B2(n_664), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_684), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_702), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_681), .A2(n_670), .B1(n_676), .B2(n_674), .C(n_668), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_684), .A2(n_288), .B1(n_293), .B2(n_302), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_699), .A2(n_302), .B(n_288), .C(n_293), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_689), .A2(n_288), .B1(n_293), .B2(n_302), .Y(n_721) );
OAI221xp5_ASAP7_75t_SL g722 ( .A1(n_695), .A2(n_293), .B1(n_302), .B2(n_685), .C(n_694), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_686), .Y(n_723) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_701), .B(n_698), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_685), .A2(n_700), .B1(n_695), .B2(n_696), .C(n_703), .Y(n_725) );
AOI211xp5_ASAP7_75t_L g726 ( .A1(n_722), .A2(n_710), .B(n_707), .C(n_714), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_713), .A2(n_725), .B1(n_709), .B2(n_718), .C(n_712), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_720), .B(n_721), .C(n_723), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_705), .B(n_706), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_708), .B(n_715), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_730), .B(n_711), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_729), .Y(n_732) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_727), .B(n_724), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_732), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_733), .A2(n_726), .B1(n_716), .B2(n_705), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_734), .Y(n_736) );
OR2x2_ASAP7_75t_SL g737 ( .A(n_735), .B(n_731), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_736), .A2(n_704), .B1(n_717), .B2(n_719), .C1(n_728), .C2(n_737), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_704), .B(n_735), .Y(n_739) );
endmodule