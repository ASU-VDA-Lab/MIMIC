module real_aes_8509_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_1), .A2(n_156), .B(n_159), .C(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_2), .A2(n_185), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g485 ( .A(n_3), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_4), .B(n_215), .Y(n_214) );
AOI21xp33_ASAP7_75t_L g468 ( .A1(n_5), .A2(n_185), .B(n_469), .Y(n_468) );
AND2x6_ASAP7_75t_L g156 ( .A(n_6), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g252 ( .A(n_7), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_42), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_8), .B(n_42), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_9), .A2(n_184), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_10), .B(n_168), .Y(n_241) );
INVx1_ASAP7_75t_L g473 ( .A(n_11), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_12), .B(n_209), .Y(n_508) );
INVx1_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
INVx1_ASAP7_75t_L g520 ( .A(n_14), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_15), .A2(n_78), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_15), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_16), .A2(n_193), .B(n_274), .C(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_17), .B(n_215), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_18), .B(n_451), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_19), .B(n_185), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_20), .B(n_199), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_21), .A2(n_209), .B(n_260), .C(n_262), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_22), .B(n_215), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_23), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_24), .A2(n_195), .B(n_276), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_25), .B(n_168), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_26), .Y(n_150) );
INVx1_ASAP7_75t_L g222 ( .A(n_27), .Y(n_222) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_28), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_29), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_30), .B(n_168), .Y(n_486) );
INVx1_ASAP7_75t_L g191 ( .A(n_31), .Y(n_191) );
INVx1_ASAP7_75t_L g463 ( .A(n_32), .Y(n_463) );
INVx2_ASAP7_75t_L g154 ( .A(n_33), .Y(n_154) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_34), .A2(n_127), .B1(n_130), .B2(n_723), .C1(n_724), .C2(n_726), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_35), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_36), .A2(n_209), .B(n_210), .C(n_212), .Y(n_208) );
INVxp67_ASAP7_75t_L g194 ( .A(n_37), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g207 ( .A(n_38), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_39), .A2(n_159), .B(n_221), .C(n_225), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_40), .A2(n_156), .B(n_159), .C(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_41), .A2(n_102), .B1(n_111), .B2(n_739), .Y(n_101) );
INVx1_ASAP7_75t_L g462 ( .A(n_43), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_44), .A2(n_170), .B(n_250), .C(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_45), .B(n_168), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_46), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_47), .Y(n_187) );
INVx1_ASAP7_75t_L g258 ( .A(n_48), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_49), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_50), .A2(n_60), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_50), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_51), .B(n_185), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_52), .A2(n_159), .B1(n_262), .B2(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_53), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_54), .Y(n_482) );
CKINVDCx14_ASAP7_75t_R g248 ( .A(n_55), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_56), .A2(n_212), .B(n_250), .C(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_57), .Y(n_125) );
INVx1_ASAP7_75t_L g470 ( .A(n_58), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_59), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_60), .Y(n_736) );
INVx1_ASAP7_75t_L g157 ( .A(n_61), .Y(n_157) );
INVx1_ASAP7_75t_L g147 ( .A(n_62), .Y(n_147) );
INVx1_ASAP7_75t_SL g211 ( .A(n_63), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_65), .B(n_215), .Y(n_264) );
INVx1_ASAP7_75t_L g163 ( .A(n_66), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_SL g450 ( .A1(n_67), .A2(n_212), .B(n_451), .C(n_452), .Y(n_450) );
INVxp67_ASAP7_75t_L g453 ( .A(n_68), .Y(n_453) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_70), .A2(n_185), .B(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_71), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_72), .A2(n_185), .B(n_271), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_73), .Y(n_466) );
INVx1_ASAP7_75t_L g526 ( .A(n_74), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_75), .A2(n_184), .B(n_186), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_76), .Y(n_219) );
INVx1_ASAP7_75t_L g272 ( .A(n_77), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_78), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_79), .A2(n_156), .B(n_159), .C(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_80), .A2(n_185), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g275 ( .A(n_81), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_82), .B(n_192), .Y(n_497) );
INVx2_ASAP7_75t_L g145 ( .A(n_83), .Y(n_145) );
INVx1_ASAP7_75t_L g240 ( .A(n_84), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_85), .B(n_451), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_86), .A2(n_156), .B(n_159), .C(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g438 ( .A(n_87), .B(n_122), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_88), .A2(n_159), .B(n_162), .C(n_172), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_89), .B(n_177), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_90), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_91), .A2(n_156), .B(n_159), .C(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_92), .Y(n_512) );
INVx1_ASAP7_75t_L g449 ( .A(n_93), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_94), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_95), .B(n_192), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_96), .B(n_143), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_97), .B(n_143), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g261 ( .A(n_99), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_100), .A2(n_185), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g740 ( .A(n_103), .Y(n_740) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g722 ( .A(n_107), .B(n_122), .Y(n_722) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_107), .B(n_121), .Y(n_728) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_126), .B1(n_729), .B2(n_731), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g730 ( .A(n_115), .Y(n_730) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_117), .A2(n_732), .B(n_737), .Y(n_731) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_125), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g738 ( .A(n_120), .Y(n_738) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g723 ( .A(n_127), .Y(n_723) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_438), .B1(n_439), .B2(n_720), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_131), .A2(n_132), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_132), .A2(n_438), .B1(n_720), .B2(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_372), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_301), .C(n_331), .D(n_352), .E(n_358), .Y(n_133) );
AOI221xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_231), .B1(n_265), .B2(n_267), .C(n_278), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_228), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_200), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_SL g352 ( .A1(n_139), .A2(n_216), .B(n_353), .C(n_356), .Y(n_352) );
AND2x2_ASAP7_75t_L g422 ( .A(n_139), .B(n_217), .Y(n_422) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_178), .Y(n_139) );
AND2x2_ASAP7_75t_L g280 ( .A(n_140), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g284 ( .A(n_140), .B(n_281), .Y(n_284) );
OR2x2_ASAP7_75t_L g310 ( .A(n_140), .B(n_217), .Y(n_310) );
AND2x2_ASAP7_75t_L g312 ( .A(n_140), .B(n_203), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_140), .B(n_202), .Y(n_330) );
INVx1_ASAP7_75t_L g363 ( .A(n_140), .Y(n_363) );
INVx2_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g230 ( .A(n_141), .Y(n_230) );
AND2x2_ASAP7_75t_L g266 ( .A(n_141), .B(n_203), .Y(n_266) );
AND2x2_ASAP7_75t_L g419 ( .A(n_141), .B(n_217), .Y(n_419) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_149), .B(n_174), .Y(n_141) );
INVx3_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_142), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_142), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g499 ( .A(n_142), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_143), .A2(n_447), .B(n_454), .Y(n_446) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_145), .B(n_146), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_158), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_151), .A2(n_177), .B(n_219), .C(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_151), .A2(n_237), .B(n_238), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_151), .A2(n_173), .B1(n_460), .B2(n_464), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_151), .A2(n_482), .B(n_483), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_151), .A2(n_526), .B(n_527), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
AND2x4_ASAP7_75t_L g185 ( .A(n_152), .B(n_156), .Y(n_185) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
INVx1_ASAP7_75t_L g263 ( .A(n_154), .Y(n_263) );
INVx1_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
INVx3_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx1_ASAP7_75t_L g451 ( .A(n_155), .Y(n_451) );
INVx4_ASAP7_75t_SL g173 ( .A(n_156), .Y(n_173) );
BUFx3_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
INVx5_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx3_ASAP7_75t_L g171 ( .A(n_160), .Y(n_171) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_167), .C(n_169), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_164), .A2(n_169), .B(n_240), .C(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_165), .A2(n_166), .B1(n_462), .B2(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx4_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
INVx2_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_169), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_169), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g276 ( .A(n_171), .Y(n_276) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g186 ( .A1(n_173), .A2(n_187), .B(n_188), .C(n_189), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_188), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_173), .A2(n_188), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_173), .A2(n_188), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_173), .A2(n_188), .B(n_272), .C(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_173), .A2(n_188), .B(n_449), .C(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_173), .A2(n_188), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_173), .A2(n_188), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_176), .A2(n_504), .B(n_511), .Y(n_503) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_177), .A2(n_246), .B(n_253), .Y(n_245) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_177), .A2(n_515), .B(n_521), .Y(n_514) );
AND2x2_ASAP7_75t_L g300 ( .A(n_178), .B(n_201), .Y(n_300) );
OR2x2_ASAP7_75t_L g304 ( .A(n_178), .B(n_217), .Y(n_304) );
AND2x2_ASAP7_75t_L g329 ( .A(n_178), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g376 ( .A(n_178), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_178), .B(n_338), .Y(n_424) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_197), .Y(n_178) );
INVx1_ASAP7_75t_L g282 ( .A(n_179), .Y(n_282) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_179), .A2(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_SL g493 ( .A1(n_180), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_181), .A2(n_459), .B(n_465), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_181), .B(n_466), .Y(n_465) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_181), .A2(n_481), .B(n_488), .Y(n_480) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_183), .A2(n_198), .B(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_190), .B(n_196), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B1(n_194), .B2(n_195), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_192), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_193), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_193), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_193), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_195), .B(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_195), .B(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_195), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI322xp33_ASAP7_75t_L g425 ( .A1(n_200), .A2(n_361), .A3(n_384), .B1(n_405), .B2(n_426), .C1(n_428), .C2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_201), .B(n_281), .Y(n_428) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
AND2x2_ASAP7_75t_L g229 ( .A(n_202), .B(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g297 ( .A(n_202), .B(n_217), .Y(n_297) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g338 ( .A(n_203), .B(n_217), .Y(n_338) );
AND2x2_ASAP7_75t_L g382 ( .A(n_203), .B(n_216), .Y(n_382) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_214), .Y(n_203) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_204), .A2(n_256), .B(n_264), .Y(n_255) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_204), .A2(n_270), .B(n_277), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_209), .B(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_213), .Y(n_509) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_215), .A2(n_468), .B(n_474), .Y(n_467) );
AND2x2_ASAP7_75t_L g265 ( .A(n_216), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g283 ( .A(n_216), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_216), .B(n_312), .Y(n_436) );
INVx3_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g228 ( .A(n_217), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_217), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g350 ( .A(n_217), .B(n_281), .Y(n_350) );
AND2x2_ASAP7_75t_L g377 ( .A(n_217), .B(n_312), .Y(n_377) );
OR2x2_ASAP7_75t_L g433 ( .A(n_217), .B(n_284), .Y(n_433) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_226), .Y(n_217) );
INVx1_ASAP7_75t_SL g319 ( .A(n_228), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_229), .B(n_350), .Y(n_351) );
AND2x2_ASAP7_75t_L g385 ( .A(n_229), .B(n_375), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_229), .B(n_308), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_229), .B(n_430), .Y(n_429) );
OAI31xp33_ASAP7_75t_L g403 ( .A1(n_231), .A2(n_265), .A3(n_404), .B(n_406), .Y(n_403) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_244), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_232), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g386 ( .A(n_232), .B(n_321), .Y(n_386) );
OR2x2_ASAP7_75t_L g393 ( .A(n_232), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g405 ( .A(n_232), .B(n_294), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g339 ( .A(n_233), .B(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g267 ( .A(n_234), .B(n_268), .Y(n_267) );
INVx4_ASAP7_75t_L g288 ( .A(n_234), .Y(n_288) );
AND2x2_ASAP7_75t_L g325 ( .A(n_234), .B(n_269), .Y(n_325) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_242), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_235), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_235), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_235), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g324 ( .A(n_244), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g394 ( .A(n_244), .Y(n_394) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_245), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_255), .Y(n_294) );
INVx2_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
AND2x2_ASAP7_75t_L g328 ( .A(n_245), .B(n_255), .Y(n_328) );
AND2x2_ASAP7_75t_L g335 ( .A(n_245), .B(n_291), .Y(n_335) );
BUFx3_ASAP7_75t_L g345 ( .A(n_245), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_245), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g290 ( .A(n_254), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_254), .B(n_288), .Y(n_298) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g268 ( .A(n_255), .B(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
INVx2_ASAP7_75t_L g487 ( .A(n_262), .Y(n_487) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_SL g305 ( .A(n_266), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_266), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_266), .B(n_375), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_267), .B(n_345), .Y(n_398) );
INVx1_ASAP7_75t_SL g432 ( .A(n_267), .Y(n_432) );
INVx1_ASAP7_75t_SL g340 ( .A(n_268), .Y(n_340) );
INVx1_ASAP7_75t_SL g291 ( .A(n_269), .Y(n_291) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_269), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_269), .B(n_288), .Y(n_313) );
AND2x2_ASAP7_75t_L g327 ( .A(n_269), .B(n_288), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_269), .B(n_317), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_283), .B(n_285), .C(n_296), .Y(n_278) );
AOI31xp33_ASAP7_75t_L g395 ( .A1(n_279), .A2(n_396), .A3(n_397), .B(n_398), .Y(n_395) );
AND2x2_ASAP7_75t_L g368 ( .A(n_280), .B(n_297), .Y(n_368) );
BUFx3_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_281), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g344 ( .A(n_281), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_281), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g299 ( .A(n_284), .Y(n_299) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_284), .A2(n_409), .B1(n_412), .B2(n_413), .C1(n_414), .C2(n_415), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_292), .Y(n_285) );
INVx1_ASAP7_75t_L g414 ( .A(n_286), .Y(n_414) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_288), .B(n_291), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_288), .B(n_314), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_288), .B(n_289), .Y(n_384) );
INVx1_ASAP7_75t_L g435 ( .A(n_288), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_289), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g437 ( .A(n_289), .Y(n_437) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
AOI32xp33_ASAP7_75t_L g296 ( .A1(n_292), .A2(n_297), .A3(n_298), .B1(n_299), .B2(n_300), .Y(n_296) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_294), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g371 ( .A(n_294), .Y(n_371) );
OR2x2_ASAP7_75t_L g412 ( .A(n_294), .B(n_313), .Y(n_412) );
INVx1_ASAP7_75t_L g348 ( .A(n_295), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_297), .B(n_308), .Y(n_333) );
INVx3_ASAP7_75t_L g342 ( .A(n_297), .Y(n_342) );
AOI322xp5_ASAP7_75t_L g358 ( .A1(n_297), .A2(n_342), .A3(n_359), .B1(n_361), .B2(n_364), .C1(n_368), .C2(n_369), .Y(n_358) );
AND2x2_ASAP7_75t_L g334 ( .A(n_298), .B(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
A2O1A1O1Ixp25_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_306), .C(n_314), .D(n_315), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_302), .B(n_345), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_304), .A2(n_316), .B1(n_319), .B2(n_320), .C(n_323), .Y(n_315) );
INVx1_ASAP7_75t_SL g430 ( .A(n_304), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B(n_313), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_308), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_310), .A2(n_394), .B1(n_401), .B2(n_402), .C(n_403), .Y(n_400) );
OAI222xp33_ASAP7_75t_L g431 ( .A1(n_311), .A2(n_432), .B1(n_433), .B2(n_434), .C1(n_436), .C2(n_437), .Y(n_431) );
AND2x2_ASAP7_75t_L g389 ( .A(n_312), .B(n_375), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_312), .A2(n_327), .B(n_374), .Y(n_401) );
INVx1_ASAP7_75t_L g415 ( .A(n_312), .Y(n_415) );
INVx2_ASAP7_75t_SL g318 ( .A(n_313), .Y(n_318) );
AND2x2_ASAP7_75t_L g321 ( .A(n_314), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_SL g355 ( .A(n_317), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_317), .B(n_327), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_318), .B(n_328), .Y(n_357) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI21xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_326), .B(n_329), .Y(n_323) );
INVx1_ASAP7_75t_SL g341 ( .A(n_325), .Y(n_341) );
AND2x2_ASAP7_75t_L g388 ( .A(n_325), .B(n_371), .Y(n_388) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g427 ( .A(n_327), .B(n_345), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_328), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g413 ( .A(n_329), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B1(n_336), .B2(n_343), .C(n_346), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B1(n_341), .B2(n_342), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_340), .A2(n_347), .B1(n_349), .B2(n_351), .Y(n_346) );
OR2x2_ASAP7_75t_L g417 ( .A(n_341), .B(n_345), .Y(n_417) );
OR2x2_ASAP7_75t_L g420 ( .A(n_341), .B(n_355), .Y(n_420) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_362), .A2(n_417), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND3xp33_ASAP7_75t_SL g372 ( .A(n_373), .B(n_387), .C(n_399), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_380), .B2(n_383), .C1(n_385), .C2(n_386), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_375), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_387) );
INVx1_ASAP7_75t_L g402 ( .A(n_388), .Y(n_402) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_L g421 ( .A1(n_392), .A2(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
NOR5xp2_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .C(n_416), .D(n_425), .E(n_431), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g725 ( .A(n_439), .Y(n_725) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_440), .B(n_657), .Y(n_439) );
NOR4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_587), .C(n_618), .D(n_637), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_545), .C(n_560), .D(n_578), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_490), .B1(n_522), .B2(n_533), .C1(n_538), .C2(n_540), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_475), .Y(n_443) );
INVx1_ASAP7_75t_L g601 ( .A(n_444), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .Y(n_444) );
AND2x2_ASAP7_75t_L g476 ( .A(n_445), .B(n_467), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_445), .B(n_479), .Y(n_630) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g537 ( .A(n_446), .B(n_457), .Y(n_537) );
AND2x2_ASAP7_75t_L g546 ( .A(n_446), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g572 ( .A(n_446), .Y(n_572) );
AND2x2_ASAP7_75t_L g593 ( .A(n_446), .B(n_457), .Y(n_593) );
BUFx2_ASAP7_75t_L g616 ( .A(n_446), .Y(n_616) );
AND2x2_ASAP7_75t_L g640 ( .A(n_446), .B(n_458), .Y(n_640) );
AND2x2_ASAP7_75t_L g704 ( .A(n_446), .B(n_467), .Y(n_704) );
AND2x2_ASAP7_75t_L g605 ( .A(n_455), .B(n_536), .Y(n_605) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_456), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
OR2x2_ASAP7_75t_L g565 ( .A(n_457), .B(n_480), .Y(n_565) );
AND2x2_ASAP7_75t_L g577 ( .A(n_457), .B(n_536), .Y(n_577) );
BUFx2_ASAP7_75t_L g709 ( .A(n_457), .Y(n_709) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g478 ( .A(n_458), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g559 ( .A(n_458), .B(n_480), .Y(n_559) );
AND2x2_ASAP7_75t_L g612 ( .A(n_458), .B(n_467), .Y(n_612) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_458), .Y(n_648) );
AND2x2_ASAP7_75t_L g535 ( .A(n_467), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g547 ( .A(n_467), .Y(n_547) );
INVx2_ASAP7_75t_L g558 ( .A(n_467), .Y(n_558) );
BUFx2_ASAP7_75t_L g582 ( .A(n_467), .Y(n_582) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_467), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AOI332xp33_ASAP7_75t_L g560 ( .A1(n_476), .A2(n_561), .A3(n_565), .B1(n_566), .B2(n_570), .B3(n_573), .C1(n_574), .C2(n_576), .Y(n_560) );
NAND2x1_ASAP7_75t_L g645 ( .A(n_476), .B(n_536), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_476), .B(n_550), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_SL g578 ( .A1(n_477), .A2(n_579), .B(n_582), .C(n_583), .Y(n_578) );
AND2x2_ASAP7_75t_L g717 ( .A(n_477), .B(n_558), .Y(n_717) );
INVx3_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g614 ( .A(n_478), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g619 ( .A(n_478), .B(n_616), .Y(n_619) );
INVx1_ASAP7_75t_L g550 ( .A(n_479), .Y(n_550) );
AND2x2_ASAP7_75t_L g653 ( .A(n_479), .B(n_612), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_479), .B(n_593), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_479), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_479), .B(n_571), .Y(n_679) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g536 ( .A(n_480), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g718 ( .A1(n_490), .A2(n_639), .A3(n_646), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
AND2x2_ASAP7_75t_L g522 ( .A(n_491), .B(n_523), .Y(n_522) );
NAND2x1_ASAP7_75t_SL g541 ( .A(n_491), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_491), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_491), .B(n_544), .Y(n_633) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_492), .A2(n_546), .B(n_548), .C(n_551), .Y(n_545) );
OR2x2_ASAP7_75t_L g562 ( .A(n_492), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g575 ( .A(n_492), .Y(n_575) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_524), .Y(n_581) );
INVx2_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
AND2x2_ASAP7_75t_L g610 ( .A(n_492), .B(n_564), .Y(n_610) );
AND2x2_ASAP7_75t_L g642 ( .A(n_492), .B(n_600), .Y(n_642) );
AND2x2_ASAP7_75t_L g646 ( .A(n_492), .B(n_569), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_492), .B(n_501), .Y(n_651) );
AND2x2_ASAP7_75t_L g685 ( .A(n_492), .B(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_492), .B(n_588), .Y(n_719) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_501), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g627 ( .A(n_501), .Y(n_627) );
AND2x2_ASAP7_75t_L g689 ( .A(n_501), .B(n_610), .Y(n_689) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
OR2x2_ASAP7_75t_L g543 ( .A(n_502), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g553 ( .A(n_502), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_502), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g661 ( .A(n_502), .Y(n_661) );
AND2x2_ASAP7_75t_L g678 ( .A(n_502), .B(n_524), .Y(n_678) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g569 ( .A(n_503), .B(n_513), .Y(n_569) );
AND2x2_ASAP7_75t_L g598 ( .A(n_503), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g609 ( .A(n_503), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_503), .B(n_564), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g523 ( .A(n_514), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g544 ( .A(n_514), .Y(n_544) );
AND2x2_ASAP7_75t_L g600 ( .A(n_514), .B(n_564), .Y(n_600) );
INVx1_ASAP7_75t_L g702 ( .A(n_522), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_523), .Y(n_706) );
INVx2_ASAP7_75t_L g564 ( .A(n_524), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_535), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_535), .B(n_640), .Y(n_698) );
OR2x2_ASAP7_75t_L g539 ( .A(n_536), .B(n_537), .Y(n_539) );
INVx1_ASAP7_75t_SL g591 ( .A(n_536), .Y(n_591) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_542), .A2(n_595), .B1(n_597), .B2(n_601), .C(n_602), .Y(n_594) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g622 ( .A(n_543), .B(n_586), .Y(n_622) );
INVx2_ASAP7_75t_L g554 ( .A(n_544), .Y(n_554) );
INVx1_ASAP7_75t_L g580 ( .A(n_544), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_544), .B(n_564), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_544), .B(n_567), .Y(n_674) );
INVx1_ASAP7_75t_L g682 ( .A(n_544), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_546), .B(n_550), .Y(n_596) );
AND2x4_ASAP7_75t_L g571 ( .A(n_547), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g684 ( .A(n_550), .B(n_640), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_553), .B(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_L g692 ( .A(n_554), .Y(n_692) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g592 ( .A(n_558), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g664 ( .A(n_558), .B(n_640), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_558), .B(n_577), .Y(n_670) );
AOI322xp5_ASAP7_75t_L g624 ( .A1(n_559), .A2(n_593), .A3(n_600), .B1(n_625), .B2(n_628), .C1(n_629), .C2(n_631), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_559), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g690 ( .A(n_562), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
INVx2_ASAP7_75t_L g567 ( .A(n_564), .Y(n_567) );
INVx1_ASAP7_75t_L g626 ( .A(n_564), .Y(n_626) );
CKINVDCx16_ASAP7_75t_R g573 ( .A(n_565), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g662 ( .A(n_567), .B(n_575), .Y(n_662) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g574 ( .A(n_569), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g617 ( .A(n_569), .B(n_610), .Y(n_617) );
AND2x2_ASAP7_75t_L g621 ( .A(n_569), .B(n_581), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_570), .A2(n_632), .B(n_634), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_570), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_701) );
INVx3_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g576 ( .A(n_571), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_571), .B(n_591), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_573), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g713 ( .A(n_580), .Y(n_713) );
INVx4_ASAP7_75t_L g586 ( .A(n_581), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_581), .B(n_608), .Y(n_656) );
INVx1_ASAP7_75t_SL g668 ( .A(n_582), .Y(n_668) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_586), .B(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_594), .C(n_611), .Y(n_587) );
OAI221xp5_ASAP7_75t_SL g707 ( .A1(n_589), .A2(n_627), .B1(n_706), .B2(n_708), .C(n_710), .Y(n_707) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_591), .B(n_704), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g683 ( .A1(n_592), .A2(n_669), .A3(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g623 ( .A(n_593), .Y(n_623) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g673 ( .A(n_598), .Y(n_673) );
AND2x2_ASAP7_75t_L g686 ( .A(n_600), .B(n_609), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_606), .Y(n_602) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_610), .B(n_713), .Y(n_712) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_620), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_619), .A2(n_688), .B(n_690), .C(n_693), .Y(n_687) );
CKINVDCx16_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_622), .B(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g649 ( .A(n_630), .Y(n_649) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_633), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g677 ( .A(n_633), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B(n_643), .C(n_652), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_641), .A2(n_651), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_714) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B1(n_647), .B2(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_SL g715 ( .A(n_654), .Y(n_715) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g657 ( .A(n_658), .B(n_687), .C(n_707), .D(n_714), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_663), .B(n_665), .C(n_683), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B(n_671), .C(n_675), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g694 ( .A(n_672), .Y(n_694) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
OR2x2_ASAP7_75t_L g705 ( .A(n_673), .B(n_706), .Y(n_705) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B(n_680), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_704), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
endmodule