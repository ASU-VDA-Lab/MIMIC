module fake_jpeg_24895_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_2),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_52),
.B1(n_47),
.B2(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_61),
.B1(n_81),
.B2(n_84),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_18),
.B1(n_37),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_18),
.B1(n_37),
.B2(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_18),
.B1(n_30),
.B2(n_33),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_28),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_83),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_72),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_29),
.B1(n_25),
.B2(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_21),
.C(n_39),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_29),
.B1(n_34),
.B2(n_39),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_34),
.B1(n_26),
.B2(n_27),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_26),
.B1(n_38),
.B2(n_85),
.Y(n_125)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_41),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_70),
.C(n_41),
.Y(n_126)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_82),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_1),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_20),
.B(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_21),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_115),
.Y(n_131)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx5_ASAP7_75t_SL g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_12),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_1),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_125),
.A2(n_137),
.B1(n_159),
.B2(n_98),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_126),
.B(n_87),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_129),
.B1(n_151),
.B2(n_157),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_55),
.B1(n_76),
.B2(n_73),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_50),
.B1(n_72),
.B2(n_67),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_130),
.A2(n_141),
.B1(n_153),
.B2(n_126),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_70),
.B(n_50),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_117),
.B(n_104),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_138),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_107),
.B1(n_109),
.B2(n_122),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_48),
.B1(n_66),
.B2(n_43),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_103),
.A2(n_48),
.B1(n_40),
.B2(n_20),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_40),
.C(n_20),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_145),
.B(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_112),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_89),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_94),
.A2(n_40),
.B1(n_2),
.B2(n_1),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_40),
.C(n_2),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_123),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_92),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_9),
.C(n_3),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_93),
.B(n_4),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_165),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_168),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_90),
.Y(n_165)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_171),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_127),
.B(n_143),
.Y(n_208)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_123),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_93),
.B1(n_114),
.B2(n_99),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_108),
.B1(n_97),
.B2(n_113),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_185),
.B1(n_194),
.B2(n_143),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_135),
.A2(n_87),
.B(n_91),
.C(n_116),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_7),
.B(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_107),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_145),
.C(n_131),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_156),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_139),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_219),
.Y(n_246)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_151),
.A3(n_139),
.B1(n_149),
.B2(n_142),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_207),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_142),
.C(n_127),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_218),
.B1(n_189),
.B2(n_163),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_215),
.B1(n_184),
.B2(n_175),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_122),
.C(n_148),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_221),
.Y(n_245)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_214),
.Y(n_233)
);

AO21x2_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_148),
.B(n_8),
.Y(n_215)
);

OA21x2_ASAP7_75t_SL g219 ( 
.A1(n_160),
.A2(n_7),
.B(n_9),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_12),
.C(n_13),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_190),
.B1(n_171),
.B2(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_232),
.B1(n_215),
.B2(n_199),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_227),
.B(n_229),
.Y(n_268)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_234),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_189),
.B1(n_175),
.B2(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_215),
.Y(n_255)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_198),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_160),
.B1(n_181),
.B2(n_172),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_213),
.C(n_207),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_258),
.C(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_248),
.B1(n_217),
.B2(n_204),
.Y(n_279)
);

AOI21x1_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_215),
.B(n_211),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_206),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_195),
.C(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.C(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_196),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_197),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_242),
.B1(n_226),
.B2(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_217),
.B1(n_245),
.B2(n_244),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_285),
.B(n_253),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_167),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_221),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_281),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_210),
.C(n_200),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_256),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_273),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_262),
.B1(n_265),
.B2(n_228),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_283),
.B1(n_279),
.B2(n_280),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_295),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_263),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_300),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_255),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_298),
.B(n_275),
.Y(n_305)
);

AOI321xp33_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_266),
.A3(n_257),
.B1(n_261),
.B2(n_249),
.C(n_246),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_277),
.C(n_281),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.C(n_309),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_277),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_290),
.B1(n_288),
.B2(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_201),
.C(n_177),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_163),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_294),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_316),
.C(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_298),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_314),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_304),
.B1(n_303),
.B2(n_174),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_180),
.C(n_14),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_312),
.Y(n_326)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_311),
.B(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_326),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_324),
.B1(n_325),
.B2(n_317),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_13),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_16),
.B(n_106),
.Y(n_333)
);


endmodule