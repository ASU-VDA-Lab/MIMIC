module fake_netlist_6_1390_n_106 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_106);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_106;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

AOI211xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_20),
.B(n_32),
.C(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2x1p5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NAND2x1p5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_45),
.B(n_42),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_30),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_44),
.B(n_45),
.C(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

OAI21x1_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_59),
.B(n_60),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

OAI21x1_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_52),
.B(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_54),
.B(n_51),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2x1p5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_62),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_43),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_74),
.Y(n_86)
);

AOI222xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_72),
.B1(n_38),
.B2(n_50),
.C1(n_67),
.C2(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_67),
.B1(n_54),
.B2(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

OAI211xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_83),
.B(n_87),
.C(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_82),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_96),
.C(n_95),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

AND3x4_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.C(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_92),
.B1(n_67),
.B2(n_1),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_92),
.B1(n_6),
.B2(n_63),
.C(n_16),
.Y(n_106)
);


endmodule