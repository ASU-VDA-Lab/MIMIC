module fake_jpeg_19241_n_291 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_22),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_13),
.B(n_25),
.C(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_13),
.B1(n_24),
.B2(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_43),
.B1(n_33),
.B2(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_13),
.B1(n_24),
.B2(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_33),
.B1(n_36),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_67),
.B1(n_48),
.B2(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_88)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_61),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_36),
.B1(n_30),
.B2(n_13),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_48),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_42),
.B(n_19),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_74),
.B1(n_85),
.B2(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_75),
.B1(n_81),
.B2(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_48),
.B1(n_45),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_53),
.B1(n_56),
.B2(n_50),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_38),
.B(n_19),
.C(n_27),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_40),
.C(n_35),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_34),
.C(n_55),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_42),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_46),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_35),
.B1(n_34),
.B2(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_67),
.B1(n_51),
.B2(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_110),
.B1(n_72),
.B2(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_62),
.B1(n_54),
.B2(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_103),
.B1(n_95),
.B2(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_79),
.B1(n_70),
.B2(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_32),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_105),
.B(n_80),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_62),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_87),
.C(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_25),
.B1(n_17),
.B2(n_16),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_79),
.B(n_85),
.C(n_88),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_92),
.B1(n_19),
.B2(n_69),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_80),
.B(n_88),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_81),
.B(n_85),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_119),
.C(n_123),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_23),
.B(n_17),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_55),
.C(n_57),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_76),
.B1(n_90),
.B2(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_76),
.B1(n_72),
.B2(n_77),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_90),
.C(n_73),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_69),
.Y(n_124)
);

XNOR2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_19),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_92),
.B1(n_16),
.B2(n_15),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_83),
.B1(n_73),
.B2(n_23),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_69),
.C(n_26),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_69),
.B1(n_19),
.B2(n_16),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_109),
.B1(n_104),
.B2(n_99),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_105),
.CI(n_97),
.CON(n_140),
.SN(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_128),
.B1(n_113),
.B2(n_117),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_150),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_91),
.C(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_159),
.C(n_160),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_134),
.B2(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_16),
.C(n_26),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_26),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_137),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_124),
.B(n_118),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_182),
.B(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_120),
.B1(n_113),
.B2(n_122),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_113),
.B1(n_116),
.B2(n_130),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_113),
.B1(n_131),
.B2(n_112),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_112),
.B1(n_132),
.B2(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_132),
.C(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_177),
.C(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_126),
.C(n_16),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_7),
.B(n_12),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_26),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_19),
.C(n_1),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_19),
.B(n_6),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_6),
.B(n_10),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_198),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_163),
.B1(n_179),
.B2(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_159),
.C(n_140),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_164),
.C(n_7),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_165),
.B1(n_182),
.B2(n_180),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_204),
.B(n_205),
.Y(n_224)
);

AOI32xp33_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_167),
.A3(n_173),
.B1(n_184),
.B2(n_170),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_165),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_140),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_166),
.B1(n_169),
.B2(n_155),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_192),
.B1(n_206),
.B2(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_161),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_195),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_223),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_164),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_226),
.C(n_189),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_11),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_241),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_192),
.C(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_231),
.C(n_234),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_194),
.C(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_193),
.C(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_201),
.C(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_234),
.C(n_228),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_191),
.B1(n_198),
.B2(n_7),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_216),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_252),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_223),
.B1(n_215),
.B2(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_215),
.C(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_237),
.C(n_240),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_237),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_9),
.B(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_191),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_250),
.B1(n_4),
.B2(n_9),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_243),
.B1(n_244),
.B2(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_264),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_221),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_8),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_9),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_11),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_263),
.B(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_259),
.C(n_260),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_10),
.B(n_11),
.Y(n_280)
);

AOI221xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_283)
);

OAI31xp67_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_269),
.A3(n_10),
.B(n_11),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_277),
.C(n_279),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_285),
.B(n_1),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_0),
.B(n_2),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_2),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_2),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_3),
.C(n_256),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_3),
.B(n_279),
.Y(n_291)
);


endmodule