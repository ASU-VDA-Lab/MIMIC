module fake_jpeg_28090_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_33),
.B1(n_29),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_43),
.B1(n_38),
.B2(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_29),
.B1(n_20),
.B2(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_61),
.B1(n_22),
.B2(n_35),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_95),
.B1(n_59),
.B2(n_25),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_75),
.B1(n_94),
.B2(n_26),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_81),
.B1(n_85),
.B2(n_99),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_19),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_98),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_39),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_34),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_100),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_32),
.B1(n_23),
.B2(n_30),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_40),
.C(n_34),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_91),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_35),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_48),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_56),
.B(n_34),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_24),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_40),
.B1(n_23),
.B2(n_32),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_23),
.B1(n_26),
.B2(n_24),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_59),
.B1(n_25),
.B2(n_21),
.Y(n_124)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_21),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_63),
.B1(n_93),
.B2(n_77),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_131),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_127),
.B1(n_94),
.B2(n_102),
.Y(n_136)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_63),
.A2(n_59),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_34),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_155),
.B1(n_156),
.B2(n_122),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_9),
.C(n_15),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_8),
.C(n_15),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_79),
.B1(n_95),
.B2(n_83),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_151),
.B(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_110),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_79),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_83),
.B(n_63),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_131),
.B(n_103),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_86),
.B1(n_62),
.B2(n_65),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_89),
.B1(n_99),
.B2(n_85),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_101),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_104),
.A2(n_74),
.B1(n_21),
.B2(n_84),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_124),
.B1(n_122),
.B2(n_112),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_154),
.B1(n_153),
.B2(n_148),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_178),
.B1(n_184),
.B2(n_142),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_143),
.B1(n_111),
.B2(n_157),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_130),
.B(n_132),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_179),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_110),
.B(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_110),
.B1(n_128),
.B2(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_191),
.B1(n_174),
.B2(n_180),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_129),
.B(n_126),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_149),
.B1(n_156),
.B2(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_162),
.C(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_177),
.C(n_171),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_126),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_109),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_109),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_111),
.B1(n_103),
.B2(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_109),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_194),
.A2(n_211),
.B1(n_212),
.B2(n_217),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_202),
.B1(n_219),
.B2(n_220),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_0),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_215),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_179),
.B(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_64),
.B1(n_76),
.B2(n_7),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_76),
.B1(n_7),
.B2(n_10),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_168),
.B(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_6),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_218),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_173),
.B1(n_188),
.B2(n_167),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_202),
.B1(n_209),
.B2(n_210),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_227),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_169),
.B1(n_187),
.B2(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_230),
.B1(n_234),
.B2(n_236),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_206),
.C(n_175),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_211),
.C(n_212),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_182),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_207),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_178),
.B1(n_193),
.B2(n_183),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_195),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_199),
.B(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_169),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_255),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_219),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_195),
.C(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_231),
.C(n_234),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_223),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_220),
.B(n_216),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_233),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_264),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_260),
.A2(n_237),
.B1(n_201),
.B2(n_229),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_265),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_230),
.B1(n_232),
.B2(n_208),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_273),
.B1(n_251),
.B2(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_256),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_205),
.C(n_170),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_253),
.C(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_243),
.B(n_242),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_283),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_10),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_272),
.B1(n_261),
.B2(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_15),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_264),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_280),
.C(n_269),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_275),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_2),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_280),
.B(n_11),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_12),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

AOI321xp33_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_304),
.A3(n_294),
.B1(n_299),
.B2(n_286),
.C(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_301),
.B(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_291),
.B(n_290),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_4),
.B(n_5),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_5),
.B(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_5),
.Y(n_309)
);


endmodule