module fake_jpeg_16800_n_245 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_25),
.B1(n_19),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_28),
.B1(n_19),
.B2(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_25),
.B1(n_29),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_24),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_20),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_23),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_61),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2x1_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_27),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_43),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_72),
.Y(n_115)
);

OAI22x1_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_19),
.B1(n_25),
.B2(n_20),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_80),
.B1(n_24),
.B2(n_2),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_20),
.B(n_38),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_17),
.B(n_33),
.C(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_85),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_22),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_22),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_83),
.B1(n_88),
.B2(n_91),
.Y(n_95)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_18),
.B1(n_28),
.B2(n_17),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_32),
.B1(n_24),
.B2(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_1),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_0),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_30),
.C(n_55),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_79),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_112),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_107),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_139)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_55),
.B(n_44),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_63),
.B1(n_81),
.B2(n_76),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_24),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_62),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_117),
.B(n_66),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_125),
.B1(n_134),
.B2(n_97),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_91),
.B1(n_74),
.B2(n_85),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_75),
.B1(n_70),
.B2(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_79),
.B(n_24),
.C(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_79),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_106),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_2),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_128),
.C(n_130),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_156),
.B(n_119),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_108),
.B1(n_95),
.B2(n_107),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_134),
.B1(n_133),
.B2(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_103),
.C(n_95),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_164),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_108),
.B(n_94),
.C(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_118),
.B1(n_94),
.B2(n_112),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_105),
.C(n_113),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_14),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_180),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_179),
.B1(n_182),
.B2(n_185),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_176),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_139),
.B1(n_140),
.B2(n_132),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_143),
.B1(n_106),
.B2(n_129),
.C(n_136),
.Y(n_178)
);

OA21x2_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_147),
.B(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_14),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_145),
.C(n_5),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_194),
.B(n_199),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_164),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_144),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_197),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_155),
.B1(n_158),
.B2(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_179),
.B1(n_170),
.B2(n_181),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_167),
.C(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_144),
.C(n_148),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_201),
.C(n_148),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_210),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_168),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_175),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_194),
.B1(n_171),
.B2(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_219),
.B1(n_221),
.B2(n_207),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_196),
.B(n_189),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_222),
.B(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_3),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_169),
.B1(n_191),
.B2(n_180),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_172),
.B1(n_174),
.B2(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_212),
.C(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_230),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_232)
);

NAND4xp25_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_211),
.C(n_5),
.D(n_6),
.Y(n_227)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_229),
.B1(n_7),
.B2(n_8),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_3),
.B(n_6),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_7),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_223),
.C(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_232),
.C(n_231),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_220),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_10),
.C(n_11),
.Y(n_241)
);

AO21x1_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_239),
.B(n_9),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_8),
.B(n_9),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.C(n_236),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.C(n_11),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_10),
.C(n_11),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);


endmodule