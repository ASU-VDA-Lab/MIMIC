module fake_jpeg_22954_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_35),
.B1(n_32),
.B2(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_75),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_35),
.B1(n_20),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_32),
.B1(n_36),
.B2(n_34),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_77),
.B1(n_82),
.B2(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_73),
.B1(n_79),
.B2(n_81),
.Y(n_111)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_74),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_22),
.B1(n_48),
.B2(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_36),
.B1(n_34),
.B2(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_30),
.B1(n_18),
.B2(n_19),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_88),
.Y(n_106)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_27),
.B1(n_24),
.B2(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_29),
.B1(n_2),
.B2(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_29),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_1),
.Y(n_125)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_97),
.Y(n_142)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_124),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_69),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_71),
.B1(n_84),
.B2(n_5),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_110),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_121),
.Y(n_154)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_123),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_65),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_89),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_86),
.B1(n_67),
.B2(n_61),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_128),
.A2(n_129),
.B1(n_144),
.B2(n_133),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_67),
.B1(n_53),
.B2(n_76),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_58),
.B1(n_53),
.B2(n_85),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_140),
.B1(n_122),
.B2(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_125),
.Y(n_170)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_62),
.B(n_74),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_104),
.B(n_92),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_64),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_148),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_60),
.B1(n_72),
.B2(n_63),
.Y(n_144)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_155),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_103),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_152),
.Y(n_185)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_16),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_125),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_189),
.B1(n_163),
.B2(n_136),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_165),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_99),
.B1(n_102),
.B2(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_163),
.A2(n_167),
.B1(n_188),
.B2(n_7),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_108),
.C(n_97),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_168),
.C(n_177),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_99),
.B1(n_118),
.B2(n_106),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_108),
.C(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_107),
.B(n_98),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_178),
.B(n_186),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_180),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_117),
.C(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_93),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_2),
.B(n_5),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_133),
.B(n_142),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_117),
.B1(n_114),
.B2(n_6),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_129),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_145),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_128),
.B(n_142),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_193),
.A2(n_209),
.B1(n_211),
.B2(n_218),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_198),
.B(n_187),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_203),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_149),
.B(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_181),
.B1(n_166),
.B2(n_182),
.Y(n_237)
);

AOI22x1_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_147),
.B1(n_152),
.B2(n_139),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_217),
.C(n_170),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_139),
.B1(n_155),
.B2(n_156),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_214),
.B(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_146),
.C(n_8),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_231),
.C(n_233),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_190),
.B1(n_189),
.B2(n_169),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_237),
.B1(n_211),
.B2(n_218),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_179),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_193),
.B(n_199),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_177),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_194),
.B(n_198),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_188),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_184),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_180),
.B(n_191),
.C(n_183),
.D(n_165),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_204),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_166),
.B(n_9),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_239),
.B(n_200),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_195),
.A2(n_196),
.B(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_8),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_203),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_249),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_253),
.B(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_255),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_238),
.B(n_244),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_217),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_222),
.C(n_233),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_197),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_205),
.B1(n_193),
.B2(n_225),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_193),
.B1(n_214),
.B2(n_206),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_228),
.B1(n_226),
.B2(n_242),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_262),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_209),
.B(n_202),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_226),
.C(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_256),
.C(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_255),
.B1(n_259),
.B2(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_278),
.C(n_274),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_288),
.C(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_253),
.B(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_289),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_249),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_235),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_299),
.B(n_257),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_281),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_199),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_266),
.C(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_288),
.B(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_271),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_307),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_284),
.B(n_265),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_221),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_312),
.A3(n_229),
.B1(n_243),
.B2(n_292),
.C1(n_283),
.C2(n_239),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_204),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_314),
.A3(n_308),
.B1(n_278),
.B2(n_247),
.C1(n_263),
.C2(n_209),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_286),
.A3(n_285),
.B1(n_290),
.B2(n_268),
.C1(n_232),
.C2(n_273),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_308),
.Y(n_317)
);

AOI321xp33_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_13),
.B(n_14),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_15),
.Y(n_320)
);


endmodule