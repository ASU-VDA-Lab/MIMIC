module fake_jpeg_17065_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_52),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_1),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_38),
.B1(n_45),
.B2(n_39),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_45),
.B1(n_39),
.B2(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_34),
.B1(n_41),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_36),
.B1(n_18),
.B2(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_2),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_69),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_6),
.B(n_28),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22x1_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_42),
.B1(n_17),
.B2(n_19),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_16),
.B1(n_32),
.B2(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_75),
.B1(n_12),
.B2(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_14),
.B1(n_29),
.B2(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_5),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_20),
.B1(n_9),
.B2(n_11),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_83),
.Y(n_86)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

NOR2x1p5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.C(n_82),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.C(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_77),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_90),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_93),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_86),
.Y(n_102)
);


endmodule