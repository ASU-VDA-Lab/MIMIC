module fake_jpeg_8368_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_53),
.B1(n_63),
.B2(n_68),
.Y(n_84)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_58),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_62),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_33),
.C(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_30),
.C(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_41),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_49),
.B1(n_63),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_17),
.B1(n_18),
.B2(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_80),
.B1(n_50),
.B2(n_51),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_41),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_87),
.C(n_20),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_81),
.Y(n_101)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_17),
.B1(n_38),
.B2(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_20),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_21),
.B(n_19),
.C(n_27),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_21),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_25),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_111),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_38),
.B1(n_60),
.B2(n_48),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_77),
.B1(n_83),
.B2(n_76),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_118),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_66),
.B1(n_46),
.B2(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_116),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_58),
.B(n_64),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_87),
.B(n_86),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_68),
.B1(n_34),
.B2(n_40),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_78),
.B1(n_79),
.B2(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_122),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_117),
.Y(n_131)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_50),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_50),
.B(n_24),
.C(n_27),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_24),
.B(n_27),
.C(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_57),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_83),
.B(n_73),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_108),
.B(n_105),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_133),
.B(n_138),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_134),
.B1(n_119),
.B2(n_118),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_108),
.B1(n_120),
.B2(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_85),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_92),
.B1(n_57),
.B2(n_62),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_142),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_88),
.B(n_1),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_78),
.A3(n_72),
.B1(n_43),
.B2(n_31),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_104),
.B(n_122),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_45),
.C(n_40),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_101),
.Y(n_163)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_148),
.Y(n_165)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_43),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_170),
.B(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_125),
.B(n_141),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_160),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_102),
.C(n_123),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_174),
.B(n_133),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_171),
.C(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_166),
.B1(n_124),
.B2(n_132),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_149),
.B1(n_124),
.B2(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_172),
.B1(n_147),
.B2(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_126),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_106),
.C(n_97),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_155),
.B1(n_152),
.B2(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_189),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_169),
.B(n_174),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_187),
.B(n_192),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_145),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_197),
.C(n_201),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_138),
.B(n_131),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_125),
.B(n_132),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_195),
.B(n_94),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_133),
.B(n_140),
.C(n_135),
.D(n_129),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_150),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_99),
.B(n_100),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_99),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_100),
.C(n_136),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_94),
.C(n_34),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_110),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_31),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_217),
.B1(n_222),
.B2(n_190),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_150),
.C(n_170),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_223),
.C(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_167),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_221),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_161),
.B1(n_156),
.B2(n_120),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_110),
.B(n_96),
.Y(n_216)
);

FAx1_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_188),
.CI(n_184),
.CON(n_230),
.SN(n_230)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_96),
.B1(n_70),
.B2(n_34),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_59),
.B1(n_52),
.B2(n_70),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_40),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_52),
.B1(n_34),
.B2(n_31),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_239),
.B(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_191),
.C(n_186),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_176),
.C(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_184),
.C(n_195),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.C(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_182),
.C(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_194),
.B1(n_182),
.B2(n_31),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_242),
.B1(n_222),
.B2(n_214),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_9),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_13),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_16),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_16),
.C(n_1),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_219),
.C(n_223),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_259),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_216),
.B1(n_215),
.B2(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_203),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_245),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_216),
.B(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_203),
.C(n_211),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_229),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_264),
.C(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_225),
.C(n_229),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_12),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_235),
.B1(n_219),
.B2(n_226),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_231),
.C(n_230),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_248),
.B(n_251),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_11),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_15),
.B(n_14),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_250),
.B(n_261),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_257),
.B(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_279),
.B1(n_271),
.B2(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_246),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_15),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_263),
.C(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_12),
.B(n_11),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_12),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_10),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_294),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_5),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_9),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_287),
.B1(n_283),
.B2(n_286),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_0),
.C(n_4),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_0),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_16),
.B(n_6),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_305),
.B(n_5),
.Y(n_306)
);

AOI31xp67_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_292),
.A3(n_289),
.B(n_296),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_302),
.B(n_300),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_16),
.B(n_7),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_16),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_313),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_307),
.Y(n_315)
);


endmodule