module fake_jpeg_17927_n_46 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_14),
.C(n_15),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_27),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_30),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_30),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_38),
.A3(n_27),
.B1(n_26),
.B2(n_24),
.C1(n_20),
.C2(n_17),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_20),
.Y(n_46)
);


endmodule