module fake_jpeg_29886_n_440 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_52),
.Y(n_93)
);

BUFx12f_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g142 ( 
.A(n_50),
.B(n_33),
.Y(n_142)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_67),
.Y(n_126)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_68),
.B(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g132 ( 
.A(n_75),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_38),
.B(n_12),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_92),
.B(n_12),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_108),
.Y(n_145)
);

CKINVDCx9p33_ASAP7_75t_R g105 ( 
.A(n_50),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_R g106 ( 
.A(n_47),
.B(n_29),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_23),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_121),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_39),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_29),
.Y(n_125)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_10),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_55),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_90),
.B1(n_80),
.B2(n_88),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_114),
.B1(n_83),
.B2(n_87),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_151),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_101),
.B(n_26),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_126),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_58),
.C(n_45),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_113),
.C(n_104),
.Y(n_209)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_61),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_161),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_43),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_177),
.Y(n_203)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_97),
.A2(n_43),
.B1(n_89),
.B2(n_77),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_175),
.B1(n_181),
.B2(n_132),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_43),
.B1(n_27),
.B2(n_41),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_101),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_93),
.B(n_73),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_121),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_183),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_27),
.B1(n_41),
.B2(n_25),
.Y(n_181)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_110),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_18),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_205),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_158),
.B(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_110),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_120),
.B1(n_133),
.B2(n_123),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_22),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_152),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_146),
.A3(n_157),
.B1(n_151),
.B2(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_222),
.Y(n_249)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_201),
.B1(n_179),
.B2(n_198),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_210),
.B1(n_190),
.B2(n_207),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_150),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_225),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_145),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_174),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_239),
.Y(n_258)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_171),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_169),
.C(n_118),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_155),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_170),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_209),
.C(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_241),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_199),
.C(n_194),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_203),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_261),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_256),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_234),
.B1(n_207),
.B2(n_233),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_186),
.B1(n_167),
.B2(n_153),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_259),
.B1(n_197),
.B2(n_185),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_200),
.B(n_191),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_237),
.B(n_230),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_191),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_153),
.B1(n_148),
.B2(n_172),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_200),
.C(n_169),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_154),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_216),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_273),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_220),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_278),
.B(n_246),
.Y(n_293)
);

AOI32xp33_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_239),
.A3(n_224),
.B1(n_226),
.B2(n_218),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_277),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_225),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_256),
.B(n_248),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_279),
.B(n_240),
.Y(n_300)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_283),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_226),
.B(n_238),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_204),
.B1(n_196),
.B2(n_235),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_259),
.B1(n_264),
.B2(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_254),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_287),
.B(n_26),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_253),
.A2(n_227),
.B1(n_219),
.B2(n_222),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_289),
.A2(n_204),
.B1(n_196),
.B2(n_202),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_229),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_248),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_300),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_235),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_308),
.B1(n_265),
.B2(n_266),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_261),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_166),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_249),
.C(n_261),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_252),
.C(n_244),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_313),
.C(n_278),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_254),
.B(n_260),
.Y(n_307)
);

HAxp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_284),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_267),
.A2(n_260),
.B1(n_251),
.B2(n_219),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_169),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_195),
.C(n_189),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_279),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_23),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_319),
.A2(n_327),
.B1(n_329),
.B2(n_337),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_323),
.C(n_332),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_283),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_325),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_268),
.C(n_290),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_289),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_328),
.A2(n_318),
.B1(n_311),
.B2(n_302),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_271),
.B(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_280),
.C(n_189),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_335),
.B(n_340),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_276),
.B1(n_206),
.B2(n_202),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_213),
.C(n_165),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_315),
.C(n_303),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_341),
.B1(n_184),
.B2(n_172),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_308),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_351),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_348),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_301),
.B1(n_293),
.B2(n_302),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_312),
.C(n_299),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_338),
.C(n_322),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_350),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_333),
.A2(n_296),
.B1(n_317),
.B2(n_295),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_295),
.C(n_297),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_354),
.C(n_355),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_168),
.C(n_156),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_176),
.C(n_177),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_340),
.A2(n_96),
.B(n_107),
.Y(n_356)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_109),
.B(n_34),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_357),
.B(n_334),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_361),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_144),
.C(n_148),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_324),
.C(n_122),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_160),
.B1(n_123),
.B2(n_128),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_352),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_360),
.B(n_323),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_370),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_353),
.A2(n_329),
.B(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_373),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_139),
.C(n_133),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_362),
.B(n_343),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_374),
.A2(n_377),
.B(n_381),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_349),
.C(n_347),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_380),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_348),
.A2(n_112),
.B(n_119),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_346),
.B(n_363),
.C(n_344),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_184),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_128),
.C(n_62),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_359),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_345),
.C(n_355),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_382),
.B(n_384),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_370),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_46),
.C(n_60),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_391),
.B(n_394),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_184),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_392),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_69),
.C(n_71),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_22),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_11),
.B(n_10),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_72),
.C(n_18),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_395),
.A2(n_0),
.B(n_1),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_379),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_401),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_378),
.C(n_368),
.Y(n_400)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_368),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_395),
.B1(n_386),
.B2(n_385),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_404),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_135),
.B1(n_130),
.B2(n_143),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_36),
.B1(n_41),
.B2(n_25),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_382),
.A2(n_36),
.B1(n_34),
.B2(n_18),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_406),
.B(n_407),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_9),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_36),
.C(n_34),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_409),
.Y(n_425)
);

OA21x2_ASAP7_75t_SL g409 ( 
.A1(n_400),
.A2(n_75),
.B(n_66),
.Y(n_409)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_410),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_396),
.A2(n_66),
.B(n_9),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_416),
.B(n_3),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_405),
.A2(n_41),
.B(n_25),
.Y(n_416)
);

AOI31xp67_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_0),
.A3(n_1),
.B(n_3),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_418),
.A2(n_0),
.B(n_3),
.Y(n_420)
);

AOI322xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_41),
.A3(n_25),
.B1(n_33),
.B2(n_5),
.C1(n_6),
.C2(n_0),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_419),
.B(n_420),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_421),
.Y(n_427)
);

NAND5xp2_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_33),
.C(n_41),
.D(n_25),
.E(n_7),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_424),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_4),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_417),
.B(n_4),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_408),
.C(n_415),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_425),
.C(n_5),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_413),
.C(n_411),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_429),
.A2(n_4),
.B(n_5),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_424),
.B(n_427),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_432),
.A2(n_434),
.B(n_6),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_433),
.B(n_430),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_436),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_7),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_8),
.B(n_330),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_8),
.Y(n_440)
);


endmodule