module fake_aes_5456_n_509 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_509);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_509;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_393;
wire n_135;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_40), .Y(n_72) );
BUFx6f_ASAP7_75t_L g73 ( .A(n_19), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_4), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_14), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_17), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_1), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_24), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_15), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_7), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_18), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_10), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_55), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_21), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_64), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_48), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_14), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_37), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_61), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_71), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_65), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_57), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_66), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_49), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_67), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_50), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_69), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_76), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_73), .Y(n_109) );
AND2x4_ASAP7_75t_L g110 ( .A(n_74), .B(n_0), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_74), .B(n_0), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_88), .B(n_1), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_104), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
BUFx8_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_75), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_93), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
AND2x6_ASAP7_75t_L g121 ( .A(n_84), .B(n_31), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_75), .B(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_121), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_107), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_106), .B(n_94), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_113), .B(n_87), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
BUFx10_ASAP7_75t_L g136 ( .A(n_121), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_108), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_118), .B(n_79), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_110), .B(n_79), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_117), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_105), .B(n_103), .Y(n_144) );
NOR2x1p5_ASAP7_75t_L g145 ( .A(n_112), .B(n_83), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_106), .B(n_94), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_118), .B(n_102), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_110), .B(n_83), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_114), .B(n_101), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_140), .A2(n_111), .B1(n_125), .B2(n_124), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_127), .B(n_108), .Y(n_153) );
INVx2_ASAP7_75t_SL g154 ( .A(n_143), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_151), .B(n_114), .Y(n_156) );
NAND2x1p5_ASAP7_75t_L g157 ( .A(n_130), .B(n_111), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_143), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_140), .B(n_111), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_129), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_140), .B(n_111), .Y(n_169) );
NOR2x2_ASAP7_75t_L g170 ( .A(n_148), .B(n_122), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_143), .Y(n_173) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_134), .Y(n_176) );
BUFx2_ASAP7_75t_SL g177 ( .A(n_130), .Y(n_177) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_134), .Y(n_179) );
OR2x2_ASAP7_75t_SL g180 ( .A(n_132), .B(n_122), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_142), .B(n_116), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_150), .B(n_116), .Y(n_184) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_184), .B(n_137), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_184), .B(n_137), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
O2A1O1Ixp5_ASAP7_75t_SL g191 ( .A1(n_152), .A2(n_92), .B(n_95), .C(n_96), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_161), .B(n_139), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_145), .B1(n_150), .B2(n_137), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
BUFx10_ASAP7_75t_L g197 ( .A(n_184), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_152), .A2(n_150), .B1(n_137), .B2(n_145), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_165), .A2(n_150), .B1(n_139), .B2(n_130), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_184), .B(n_139), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_164), .B(n_130), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_153), .A2(n_142), .B(n_146), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_165), .B(n_132), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_153), .A2(n_146), .B(n_144), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_184), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_160), .B(n_147), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_164), .A2(n_121), .B1(n_147), .B2(n_120), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_174), .B(n_120), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_180), .B(n_183), .Y(n_215) );
INVx4_ASAP7_75t_SL g216 ( .A(n_187), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_200), .A2(n_174), .B1(n_178), .B2(n_160), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_198), .A2(n_174), .B1(n_178), .B2(n_160), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_200), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_185), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_197), .Y(n_222) );
BUFx8_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
INVx6_ASAP7_75t_L g224 ( .A(n_197), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_198), .A2(n_174), .B1(n_178), .B2(n_160), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_197), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_200), .B(n_180), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_211), .A2(n_156), .B(n_183), .C(n_123), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_207), .A2(n_178), .B1(n_169), .B2(n_160), .Y(n_230) );
CKINVDCx9p33_ASAP7_75t_R g231 ( .A(n_204), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_205), .B(n_156), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_197), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_200), .A2(n_169), .B1(n_176), .B2(n_179), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_202), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_205), .B(n_169), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
AOI222xp33_ASAP7_75t_L g238 ( .A1(n_194), .A2(n_80), .B1(n_170), .B2(n_169), .C1(n_123), .C2(n_124), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_194), .A2(n_169), .B1(n_182), .B2(n_179), .Y(n_239) );
BUFx4f_ASAP7_75t_SL g240 ( .A(n_221), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_227), .A2(n_208), .B(n_190), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_232), .A2(n_215), .B1(n_195), .B2(n_211), .C(n_199), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_236), .B(n_214), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_229), .A2(n_215), .B1(n_214), .B2(n_125), .C(n_188), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_238), .A2(n_185), .B1(n_207), .B2(n_204), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g247 ( .A1(n_223), .A2(n_185), .B1(n_210), .B2(n_209), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_219), .A2(n_196), .B1(n_190), .B2(n_208), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_237), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_237), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_225), .A2(n_196), .B(n_208), .Y(n_252) );
BUFx4f_ASAP7_75t_SL g253 ( .A(n_223), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_196), .B1(n_213), .B2(n_210), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_218), .A2(n_213), .A3(n_192), .B(n_209), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_223), .A2(n_202), .B1(n_187), .B2(n_193), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_238), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_191), .B(n_203), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_236), .A2(n_189), .B1(n_188), .B2(n_206), .C(n_80), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_240), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_246), .A2(n_218), .B1(n_217), .B2(n_226), .Y(n_261) );
OAI33xp33_ASAP7_75t_L g262 ( .A1(n_257), .A2(n_92), .A3(n_95), .B1(n_96), .B2(n_97), .B3(n_98), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_250), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_253), .A2(n_228), .B1(n_220), .B2(n_224), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_245), .A2(n_228), .B1(n_226), .B2(n_224), .Y(n_265) );
OAI321xp33_ASAP7_75t_L g266 ( .A1(n_254), .A2(n_100), .A3(n_98), .B1(n_97), .B2(n_78), .C(n_73), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_243), .A2(n_234), .B1(n_206), .B2(n_115), .C(n_119), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_241), .A2(n_224), .B1(n_233), .B2(n_222), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_212), .B1(n_189), .B2(n_222), .C(n_233), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_252), .A2(n_191), .B(n_203), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_241), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_244), .A2(n_224), .B1(n_235), .B2(n_231), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_244), .B(n_115), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_249), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_250), .B(n_235), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_258), .A2(n_100), .B(n_119), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_248), .A2(n_162), .B(n_168), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_263), .B(n_255), .Y(n_281) );
OAI33xp33_ASAP7_75t_L g282 ( .A1(n_279), .A2(n_2), .A3(n_3), .B1(n_4), .B2(n_5), .B3(n_6), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_263), .B(n_255), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_277), .Y(n_284) );
NAND2x1_ASAP7_75t_L g285 ( .A(n_277), .B(n_249), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_262), .A2(n_259), .B1(n_91), .B2(n_99), .C(n_81), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_278), .B(n_255), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_260), .B(n_3), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_279), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_274), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_274), .B(n_258), .Y(n_293) );
AOI33xp33_ASAP7_75t_L g294 ( .A1(n_264), .A2(n_256), .A3(n_6), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_275), .B(n_242), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_273), .B(n_235), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_275), .B(n_216), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_261), .B(n_5), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_73), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_265), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_265), .A2(n_121), .B1(n_193), .B2(n_187), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_78), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_269), .A2(n_117), .B(n_193), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_272), .B(n_216), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_280), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_268), .A2(n_157), .B1(n_78), .B2(n_201), .C(n_162), .Y(n_310) );
OAI31xp33_ASAP7_75t_SL g311 ( .A1(n_267), .A2(n_216), .A3(n_10), .B(n_11), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_280), .B(n_78), .Y(n_312) );
INVx3_ASAP7_75t_SL g313 ( .A(n_298), .Y(n_313) );
OAI33xp33_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_8), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_15), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_287), .B(n_270), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_285), .Y(n_316) );
BUFx2_ASAP7_75t_SL g317 ( .A(n_298), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_12), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_281), .B(n_78), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_283), .B(n_126), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_281), .B(n_216), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_283), .B(n_126), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_300), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g327 ( .A1(n_299), .A2(n_13), .A3(n_16), .B1(n_266), .B2(n_85), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_289), .B(n_126), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_289), .B(n_16), .Y(n_329) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_282), .B(n_86), .C(n_90), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_301), .B(n_109), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_304), .A2(n_121), .B(n_157), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_281), .B(n_126), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_297), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_292), .B(n_126), .Y(n_336) );
AOI322xp5_ASAP7_75t_L g337 ( .A1(n_288), .A2(n_109), .A3(n_126), .B1(n_202), .B2(n_193), .C1(n_168), .C2(n_171), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_294), .B(n_109), .C(n_117), .Y(n_338) );
NAND5xp2_ASAP7_75t_L g339 ( .A(n_311), .B(n_157), .C(n_201), .D(n_121), .E(n_26), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_293), .B(n_20), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_297), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_293), .B(n_22), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_305), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_312), .B(n_25), .Y(n_345) );
NOR2xp33_ASAP7_75t_SL g346 ( .A(n_298), .B(n_202), .Y(n_346) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_312), .B(n_202), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_295), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_295), .B(n_121), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_307), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_296), .B(n_175), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_308), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_357), .B(n_310), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_349), .B(n_309), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_326), .B(n_302), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_313), .B(n_27), .Y(n_363) );
NOR2x1p5_ASAP7_75t_L g364 ( .A(n_316), .B(n_286), .Y(n_364) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_320), .B(n_177), .Y(n_365) );
OAI33xp33_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_117), .A3(n_175), .B1(n_172), .B2(n_171), .B3(n_181), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_320), .B(n_28), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_315), .B(n_29), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_345), .B(n_202), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_30), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_321), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_313), .B(n_34), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_322), .B(n_35), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_341), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_325), .B(n_38), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_324), .B(n_39), .Y(n_380) );
NAND2xp33_ASAP7_75t_L g381 ( .A(n_313), .B(n_202), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_324), .B(n_42), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_325), .B(n_43), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_315), .B(n_44), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_328), .Y(n_385) );
NOR2x1p5_ASAP7_75t_SL g386 ( .A(n_334), .B(n_175), .Y(n_386) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_317), .B(n_201), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_328), .B(n_45), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_319), .B(n_46), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_351), .B(n_47), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_344), .Y(n_392) );
NOR4xp25_ASAP7_75t_L g393 ( .A(n_318), .B(n_181), .C(n_172), .D(n_171), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_353), .B(n_51), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_344), .B(n_52), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_317), .B(n_53), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_333), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_348), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_347), .B(n_54), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_351), .B(n_56), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_335), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_353), .B(n_58), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_351), .B(n_59), .Y(n_404) );
OAI31xp33_ASAP7_75t_L g405 ( .A1(n_339), .A2(n_157), .A3(n_173), .B(n_154), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_347), .B(n_60), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_376), .B(n_350), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_388), .B(n_340), .Y(n_411) );
XNOR2x1_ASAP7_75t_L g412 ( .A(n_387), .B(n_338), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_360), .A2(n_314), .B1(n_330), .B2(n_346), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_397), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_381), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_327), .B(n_345), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_327), .B(n_340), .C(n_343), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_331), .B1(n_355), .B2(n_333), .C(n_343), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_402), .Y(n_424) );
NAND2xp33_ASAP7_75t_L g425 ( .A(n_363), .B(n_334), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_372), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_399), .B(n_355), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_365), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_406), .B(n_352), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_359), .B(n_335), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
XOR2x2_ASAP7_75t_L g434 ( .A(n_369), .B(n_356), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_385), .B(n_352), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_362), .B(n_358), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_374), .B(n_358), .Y(n_437) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_400), .A2(n_337), .A3(n_336), .B1(n_354), .B2(n_332), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_375), .B(n_336), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_386), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_364), .A2(n_337), .B1(n_163), .B2(n_179), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_368), .B(n_62), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_394), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_403), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_366), .B(n_63), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_405), .B(n_182), .C(n_179), .D(n_176), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_408), .A2(n_149), .B(n_135), .C(n_141), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_380), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_368), .B(n_68), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_395), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_391), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_384), .B(n_172), .C(n_181), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_389), .A2(n_163), .B1(n_176), .B2(n_182), .Y(n_455) );
AOI221x1_ASAP7_75t_L g456 ( .A1(n_384), .A2(n_135), .B1(n_149), .B2(n_141), .C(n_163), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_380), .A2(n_173), .B(n_154), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_390), .B(n_135), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_391), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_404), .B(n_135), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_382), .A2(n_163), .B1(n_176), .B2(n_182), .Y(n_462) );
XNOR2x1_ASAP7_75t_L g463 ( .A(n_382), .B(n_177), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_404), .B(n_154), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_396), .B(n_135), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_370), .A2(n_173), .B(n_141), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_367), .A2(n_135), .B1(n_141), .B2(n_149), .C(n_136), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_373), .B(n_135), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_401), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_378), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_383), .B(n_141), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_376), .B(n_149), .Y(n_472) );
AOI211xp5_ASAP7_75t_SL g473 ( .A1(n_381), .A2(n_149), .B(n_141), .C(n_136), .Y(n_473) );
NAND3x2_ASAP7_75t_L g474 ( .A(n_400), .B(n_149), .C(n_141), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_446), .B(n_447), .C(n_472), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_412), .A2(n_427), .B1(n_414), .B2(n_458), .Y(n_476) );
OA33x2_ASAP7_75t_L g477 ( .A1(n_410), .A2(n_435), .A3(n_437), .B1(n_439), .B2(n_432), .B3(n_428), .Y(n_477) );
BUFx8_ASAP7_75t_L g478 ( .A(n_450), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_415), .A2(n_452), .B1(n_422), .B2(n_470), .C(n_441), .Y(n_479) );
AOI211x1_ASAP7_75t_L g480 ( .A1(n_430), .A2(n_418), .B(n_440), .C(n_411), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_446), .A2(n_463), .B1(n_454), .B2(n_434), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
AOI31xp33_ASAP7_75t_L g484 ( .A1(n_417), .A2(n_421), .A3(n_429), .B(n_449), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_431), .Y(n_485) );
AOI322xp5_ASAP7_75t_L g486 ( .A1(n_415), .A2(n_436), .A3(n_430), .B1(n_425), .B2(n_429), .C1(n_416), .C2(n_420), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_413), .A2(n_438), .B(n_425), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_413), .A2(n_474), .B1(n_424), .B2(n_471), .Y(n_488) );
AOI21xp33_ASAP7_75t_SL g489 ( .A1(n_465), .A2(n_464), .B(n_453), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_487), .A2(n_448), .B1(n_445), .B2(n_444), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_476), .A2(n_462), .B(n_442), .C(n_455), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_478), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_480), .B(n_424), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_479), .A2(n_426), .B1(n_409), .B2(n_423), .C(n_469), .Y(n_494) );
AOI211x1_ASAP7_75t_SL g495 ( .A1(n_488), .A2(n_465), .B(n_443), .C(n_451), .Y(n_495) );
BUFx12f_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_475), .A2(n_460), .B1(n_472), .B2(n_468), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_490), .B(n_486), .C(n_481), .Y(n_498) );
NAND5xp2_ASAP7_75t_L g499 ( .A(n_494), .B(n_455), .C(n_462), .D(n_473), .E(n_484), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_492), .B(n_489), .C(n_459), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_493), .A2(n_485), .B1(n_483), .B2(n_482), .C(n_477), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_498), .B(n_495), .C(n_491), .D(n_497), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_500), .Y(n_503) );
AOI22x1_ASAP7_75t_L g504 ( .A1(n_503), .A2(n_496), .B1(n_499), .B2(n_501), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_502), .A2(n_468), .B1(n_461), .B2(n_456), .Y(n_505) );
NOR3x1_ASAP7_75t_L g506 ( .A(n_504), .B(n_457), .C(n_466), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_506), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_507), .Y(n_508) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_508), .A2(n_505), .B(n_467), .Y(n_509) );
endmodule