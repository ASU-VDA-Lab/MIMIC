module fake_aes_5938_n_739 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_739);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_739;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_553;
wire n_440;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g93 ( .A(n_65), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_19), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_39), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_91), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_21), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_40), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_10), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_34), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_18), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_50), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_53), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_54), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_6), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_75), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_69), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_12), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_85), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_28), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_1), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_12), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_86), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_88), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_1), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_72), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_112), .B(n_0), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_96), .B(n_92), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_94), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_110), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_103), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_103), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_106), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_96), .B(n_0), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx6_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_115), .B(n_2), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_100), .A2(n_41), .B(n_89), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_144), .B(n_122), .Y(n_152) );
INVx1_ASAP7_75t_SL g153 ( .A(n_133), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_144), .B(n_109), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_142), .B(n_124), .Y(n_158) );
NOR2x1p5_ASAP7_75t_L g159 ( .A(n_143), .B(n_119), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_149), .B(n_123), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_149), .B(n_127), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_150), .B(n_95), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_130), .A2(n_128), .B1(n_118), .B2(n_119), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_129), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_150), .B(n_99), .Y(n_174) );
INVxp33_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_139), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
NAND2xp33_ASAP7_75t_L g178 ( .A(n_141), .B(n_98), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_142), .A2(n_101), .B1(n_125), .B2(n_121), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_142), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_171), .B(n_142), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_174), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_171), .B(n_141), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_180), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_168), .A2(n_147), .B1(n_101), .B2(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_182), .B(n_111), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_170), .B(n_147), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_156), .B(n_148), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_160), .B(n_148), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_163), .B(n_148), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_167), .B(n_116), .Y(n_199) );
NOR2x1p5_ASAP7_75t_L g200 ( .A(n_174), .B(n_148), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_168), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_164), .B(n_134), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_151), .B(n_136), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_159), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_151), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_177), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_159), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_177), .B(n_136), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_167), .B(n_104), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_177), .B(n_131), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_167), .A2(n_131), .B1(n_137), .B2(n_105), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_166), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_172), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_179), .B(n_105), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_176), .Y(n_219) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_179), .B(n_145), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_179), .B(n_108), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_175), .A2(n_137), .B1(n_108), .B2(n_121), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_152), .B(n_158), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_183), .A2(n_137), .B1(n_113), .B2(n_125), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_154), .B(n_113), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g226 ( .A1(n_202), .A2(n_161), .B(n_154), .C(n_157), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_207), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_187), .B(n_178), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_197), .B(n_114), .Y(n_229) );
INVx1_ASAP7_75t_SL g230 ( .A(n_188), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_187), .A2(n_114), .B1(n_117), .B2(n_120), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_188), .B(n_117), .Y(n_232) );
O2A1O1Ixp5_ASAP7_75t_L g233 ( .A1(n_214), .A2(n_221), .B(n_217), .C(n_199), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_207), .B(n_157), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_223), .B(n_120), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_192), .B(n_126), .Y(n_236) );
CKINVDCx14_ASAP7_75t_R g237 ( .A(n_201), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_200), .B(n_126), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_209), .A2(n_145), .B(n_165), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_200), .B(n_135), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_222), .A2(n_135), .B(n_140), .C(n_165), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_205), .B(n_2), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_195), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_225), .A2(n_162), .B(n_173), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_209), .A2(n_145), .B(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_198), .B(n_213), .C(n_211), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_220), .A2(n_145), .B(n_161), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_220), .A2(n_173), .B(n_181), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_193), .A2(n_135), .B(n_140), .C(n_181), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_193), .A2(n_218), .B(n_219), .C(n_204), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_205), .B(n_3), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_185), .B(n_172), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_186), .B(n_135), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_218), .A2(n_185), .B(n_184), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_230), .B(n_201), .Y(n_258) );
NOR2x1_ASAP7_75t_SL g259 ( .A(n_243), .B(n_212), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_238), .B(n_210), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_255), .A2(n_219), .B(n_194), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_249), .A2(n_212), .B(n_189), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_246), .B(n_210), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_212), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_189), .B(n_194), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_238), .B(n_190), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_229), .B(n_208), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_253), .A2(n_191), .B1(n_224), .B2(n_208), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_251), .A2(n_216), .B(n_215), .Y(n_270) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_247), .A2(n_184), .A3(n_155), .B(n_206), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_227), .B(n_203), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_248), .A2(n_184), .B(n_155), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_235), .A2(n_140), .B(n_135), .C(n_155), .Y(n_274) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_245), .A2(n_216), .B(n_215), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_234), .A2(n_206), .B(n_169), .Y(n_276) );
NAND3xp33_ASAP7_75t_SL g277 ( .A(n_242), .B(n_3), .C(n_4), .Y(n_277) );
NOR3xp33_ASAP7_75t_L g278 ( .A(n_242), .B(n_4), .C(n_5), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_169), .B(n_140), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_267), .B(n_252), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_265), .A2(n_244), .B(n_240), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_275), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g283 ( .A1(n_277), .A2(n_231), .B(n_241), .C(n_236), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_261), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_271), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_273), .A2(n_256), .B(n_227), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_271), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_273), .A2(n_250), .B(n_233), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_279), .A2(n_234), .B(n_252), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_266), .B(n_235), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_258), .B(n_232), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_270), .A2(n_226), .B(n_254), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_262), .A2(n_254), .B(n_140), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_274), .A2(n_140), .A3(n_169), .B(n_7), .Y(n_295) );
OAI221xp5_ASAP7_75t_SL g296 ( .A1(n_266), .A2(n_5), .B1(n_6), .B2(n_7), .C(n_8), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_274), .A2(n_169), .B(n_45), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_267), .B(n_272), .Y(n_299) );
AO31x2_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_169), .A3(n_9), .B(n_10), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_263), .A2(n_8), .B(n_11), .C(n_13), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_292), .B(n_259), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_291), .B(n_264), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_291), .B(n_269), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_295), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_292), .B(n_263), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_296), .B(n_278), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_301), .B(n_268), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_11), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_303), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_293), .A2(n_294), .B(n_284), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_295), .B(n_13), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_280), .B(n_276), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_285), .A2(n_49), .B(n_87), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_300), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_290), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_290), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_283), .A2(n_293), .B(n_294), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_287), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_287), .Y(n_342) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_305), .B(n_296), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_337), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_316), .A2(n_283), .B(n_287), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_308), .B(n_302), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_310), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_311), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_327), .B(n_300), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_327), .B(n_297), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_342), .B(n_297), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_341), .B(n_297), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_309), .B(n_289), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_308), .B(n_313), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_309), .B(n_289), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_312), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_312), .B(n_289), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_314), .B(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_314), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_305), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_319), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_315), .B(n_298), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_320), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_307), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_331), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_319), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_331), .B(n_298), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_313), .B(n_298), .Y(n_392) );
INVx3_ASAP7_75t_L g393 ( .A(n_337), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_319), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_335), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_322), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_339), .B(n_298), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_322), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_339), .B(n_286), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_326), .B(n_281), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_318), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_322), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_334), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_307), .B(n_14), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_336), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_340), .A2(n_281), .B(n_15), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_362), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_336), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_362), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_357), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_364), .B(n_321), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_374), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_405), .B(n_325), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_402), .B(n_326), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_377), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_371), .B(n_317), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_385), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_363), .B(n_321), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_389), .B(n_338), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_378), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_405), .B(n_317), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_379), .B(n_325), .Y(n_429) );
BUFx2_ASAP7_75t_SL g430 ( .A(n_383), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_363), .B(n_321), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_385), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_384), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_359), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_349), .B(n_318), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_359), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_359), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_367), .B(n_323), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_372), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_389), .B(n_395), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_372), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_386), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_386), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_380), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_385), .B(n_330), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_370), .B(n_321), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_343), .B(n_340), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_346), .B(n_329), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_395), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_397), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_397), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_404), .B(n_407), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_370), .B(n_332), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_404), .B(n_332), .Y(n_459) );
INVx5_ASAP7_75t_L g460 ( .A(n_381), .Y(n_460) );
INVx3_ASAP7_75t_SL g461 ( .A(n_366), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_356), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_373), .B(n_338), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_373), .B(n_338), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_375), .B(n_329), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_366), .Y(n_467) );
OR2x6_ASAP7_75t_L g468 ( .A(n_407), .B(n_408), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_375), .B(n_329), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_356), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_376), .B(n_329), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_376), .B(n_330), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_408), .B(n_367), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_358), .B(n_330), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_392), .B(n_14), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_394), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_366), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_358), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_366), .B(n_16), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_396), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_360), .B(n_16), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_360), .B(n_17), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_365), .B(n_20), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_368), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_396), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_368), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_369), .B(n_22), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_399), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_369), .B(n_23), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_345), .Y(n_490) );
AND2x4_ASAP7_75t_SL g491 ( .A(n_361), .B(n_24), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_347), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_400), .B(n_25), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_347), .Y(n_494) );
NOR2xp67_ASAP7_75t_L g495 ( .A(n_344), .B(n_26), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_400), .B(n_27), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_381), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_399), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_361), .B(n_406), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_348), .B(n_29), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_413), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_473), .B(n_350), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_441), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_461), .B(n_406), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_479), .Y(n_507) );
INVx3_ASAP7_75t_SL g508 ( .A(n_430), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_424), .B(n_350), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_424), .B(n_351), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_473), .B(n_351), .Y(n_511) );
AND3x1_ASAP7_75t_L g512 ( .A(n_418), .B(n_382), .C(n_391), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_415), .B(n_354), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_411), .B(n_354), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_431), .B(n_352), .Y(n_515) );
AOI32xp33_ASAP7_75t_L g516 ( .A1(n_418), .A2(n_401), .A3(n_382), .B1(n_398), .B2(n_391), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_441), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_457), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_422), .B(n_348), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_411), .B(n_352), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_479), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_457), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_410), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_449), .A2(n_401), .B1(n_398), .B2(n_409), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_439), .B(n_353), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_412), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_493), .B(n_353), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_416), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_417), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_420), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_477), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_465), .B(n_355), .Y(n_532) );
OAI21xp33_ASAP7_75t_L g533 ( .A1(n_451), .A2(n_401), .B(n_355), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_421), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_427), .B(n_403), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_412), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_426), .Y(n_537) );
NAND2x1_ASAP7_75t_L g538 ( .A(n_468), .B(n_393), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_419), .B(n_403), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
OR3x2_ASAP7_75t_L g541 ( .A(n_429), .B(n_409), .C(n_32), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_409), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_458), .B(n_393), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_458), .B(n_393), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_393), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_467), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_469), .B(n_387), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_428), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_434), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_475), .B(n_387), .Y(n_550) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_435), .B(n_387), .C(n_344), .D(n_36), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_469), .B(n_387), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_468), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_433), .B(n_344), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_471), .B(n_344), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_446), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_431), .B(n_381), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_438), .Y(n_559) );
NOR2xp33_ASAP7_75t_SL g560 ( .A(n_493), .B(n_381), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_444), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_463), .B(n_381), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_445), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_450), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_453), .B(n_30), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_460), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_35), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_455), .B(n_37), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_456), .B(n_448), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_462), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_464), .B(n_38), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_470), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_448), .B(n_42), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_464), .B(n_43), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_450), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_481), .B(n_44), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_423), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_478), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_481), .B(n_46), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_414), .B(n_51), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_468), .B(n_55), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_414), .B(n_56), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_423), .B(n_57), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_459), .B(n_58), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_496), .B(n_60), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_484), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_459), .B(n_61), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_486), .B(n_62), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_490), .B(n_63), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_452), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_496), .B(n_64), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_432), .B(n_492), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_569), .B(n_494), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_569), .B(n_499), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_501), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_504), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_508), .B(n_432), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_518), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_522), .B(n_499), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_503), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_528), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_552), .B(n_472), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_551), .A2(n_491), .B(n_447), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_530), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_532), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_577), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_512), .B(n_425), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_548), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_559), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
NAND2x1_ASAP7_75t_L g614 ( .A(n_556), .B(n_425), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_561), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_511), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_563), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_513), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_570), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_509), .B(n_510), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_540), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_553), .B(n_425), .C(n_437), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_592), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_521), .B(n_443), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_581), .B(n_489), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_551), .A2(n_495), .B(n_487), .Y(n_626) );
NAND2x1_ASAP7_75t_SL g627 ( .A(n_556), .B(n_487), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_572), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_527), .A2(n_447), .B1(n_460), .B2(n_474), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_566), .B(n_452), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_525), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_557), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
NOR2xp33_ASAP7_75t_R g634 ( .A(n_507), .B(n_483), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_509), .B(n_485), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_575), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_510), .B(n_485), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_590), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_515), .B(n_498), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_515), .B(n_498), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_514), .B(n_440), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_578), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_577), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_523), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_520), .B(n_466), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_586), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_539), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_502), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_519), .B(n_466), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_516), .B(n_454), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_535), .Y(n_651) );
NAND2x2_ASAP7_75t_L g652 ( .A(n_538), .B(n_474), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_505), .B(n_454), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_517), .B(n_476), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_554), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_562), .B(n_437), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_595), .A2(n_573), .B(n_580), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_650), .A2(n_533), .B1(n_524), .B2(n_542), .C(n_545), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_603), .A2(n_581), .B(n_527), .Y(n_659) );
AOI321xp33_ASAP7_75t_SL g660 ( .A1(n_607), .A2(n_531), .A3(n_576), .B1(n_541), .B2(n_591), .C(n_533), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_650), .B(n_536), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_608), .A2(n_550), .B1(n_558), .B2(n_506), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_655), .B(n_526), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_620), .B(n_549), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g665 ( .A1(n_597), .A2(n_585), .A3(n_583), .B(n_567), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_601), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_647), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_594), .B(n_558), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_604), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_602), .B(n_531), .Y(n_670) );
OAI32xp33_ASAP7_75t_L g671 ( .A1(n_652), .A2(n_574), .A3(n_587), .B1(n_584), .B2(n_547), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_645), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_613), .A2(n_544), .A3(n_543), .B1(n_573), .B2(n_560), .C1(n_579), .C2(n_568), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_630), .Y(n_674) );
AO22x1_ASAP7_75t_L g675 ( .A1(n_608), .A2(n_566), .B1(n_571), .B2(n_582), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_605), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_623), .A2(n_566), .B1(n_497), .B2(n_443), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_609), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_610), .Y(n_679) );
AO32x1_ASAP7_75t_L g680 ( .A1(n_596), .A2(n_491), .A3(n_482), .B1(n_483), .B2(n_442), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_651), .B(n_568), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_631), .Y(n_682) );
AOI322xp5_ASAP7_75t_L g683 ( .A1(n_620), .A2(n_565), .A3(n_482), .B1(n_589), .B2(n_588), .C1(n_436), .C2(n_440), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_611), .Y(n_684) );
NAND2xp33_ASAP7_75t_L g685 ( .A(n_634), .B(n_460), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_618), .B(n_480), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_606), .B(n_434), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_648), .A2(n_616), .B1(n_600), .B2(n_598), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_594), .B(n_476), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_607), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_612), .Y(n_691) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_599), .A2(n_565), .A3(n_436), .B1(n_442), .B2(n_480), .C1(n_488), .C2(n_500), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_658), .A2(n_599), .B(n_593), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_671), .A2(n_615), .B1(n_617), .B2(n_619), .C(n_646), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_685), .A2(n_603), .B(n_614), .Y(n_695) );
OAI21xp33_ASAP7_75t_SL g696 ( .A1(n_659), .A2(n_627), .B(n_643), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_659), .A2(n_625), .B1(n_622), .B2(n_643), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_665), .A2(n_674), .B(n_681), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_661), .B(n_593), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_665), .A2(n_629), .B(n_628), .Y(n_700) );
OAI321xp33_ASAP7_75t_L g701 ( .A1(n_660), .A2(n_626), .A3(n_625), .B1(n_639), .B2(n_635), .C(n_653), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_662), .A2(n_626), .B1(n_635), .B2(n_639), .C(n_642), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_661), .A2(n_649), .B1(n_654), .B2(n_653), .C(n_624), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_673), .A2(n_649), .B1(n_654), .B2(n_641), .C(n_656), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_664), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_675), .A2(n_640), .B(n_637), .C(n_633), .Y(n_706) );
OAI321xp33_ASAP7_75t_L g707 ( .A1(n_660), .A2(n_621), .A3(n_632), .B1(n_638), .B2(n_636), .C(n_644), .Y(n_707) );
AOI22xp5_ASAP7_75t_SL g708 ( .A1(n_664), .A2(n_497), .B1(n_67), .B2(n_70), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_677), .A2(n_66), .B1(n_71), .B2(n_73), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_668), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_682), .A2(n_74), .B1(n_76), .B2(n_77), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_666), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_688), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_84), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_669), .B(n_90), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_667), .B(n_692), .Y(n_715) );
AOI21xp5_ASAP7_75t_SL g716 ( .A1(n_680), .A2(n_690), .B(n_678), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_680), .A2(n_686), .B(n_663), .Y(n_717) );
OAI221xp5_ASAP7_75t_SL g718 ( .A1(n_683), .A2(n_689), .B1(n_670), .B2(n_672), .C(n_676), .Y(n_718) );
AOI33xp33_ASAP7_75t_L g719 ( .A1(n_679), .A2(n_684), .A3(n_691), .B1(n_687), .B2(n_657), .B3(n_680), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_657), .B(n_658), .C(n_665), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_693), .B(n_720), .Y(n_721) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_697), .B(n_695), .Y(n_722) );
OR3x1_ASAP7_75t_L g723 ( .A(n_701), .B(n_707), .C(n_698), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_719), .B(n_718), .C(n_694), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_715), .B(n_717), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_725), .B(n_707), .C(n_696), .Y(n_726) );
NAND3xp33_ASAP7_75t_SL g727 ( .A(n_724), .B(n_706), .C(n_702), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_722), .B(n_710), .Y(n_728) );
NAND4xp25_ASAP7_75t_SL g729 ( .A(n_726), .B(n_721), .C(n_723), .D(n_716), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_727), .B(n_713), .C(n_700), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_729), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_730), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_731), .A2(n_728), .B(n_705), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_732), .B(n_712), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_733), .B(n_732), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_735), .A2(n_734), .B(n_699), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_736), .A2(n_709), .B(n_708), .Y(n_737) );
AO21x2_ASAP7_75t_L g738 ( .A1(n_737), .A2(n_711), .B(n_714), .Y(n_738) );
AOI21xp33_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_704), .B(n_703), .Y(n_739) );
endmodule