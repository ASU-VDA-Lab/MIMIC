module fake_aes_11448_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI21x1_ASAP7_75t_L g12 ( .A1(n_3), .A2(n_2), .B(n_11), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_5), .B(n_1), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_13), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR4xp25_ASAP7_75t_L g22 ( .A(n_19), .B(n_17), .C(n_14), .D(n_15), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_16), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_21), .B(n_16), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_19), .B1(n_17), .B2(n_13), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_25), .B1(n_20), .B2(n_13), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_28), .B(n_0), .Y(n_29) );
NOR2x1p5_ASAP7_75t_L g30 ( .A(n_27), .B(n_13), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_1), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_31), .B(n_4), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_12), .B1(n_18), .B2(n_6), .Y(n_33) );
NAND3xp33_ASAP7_75t_SL g34 ( .A(n_29), .B(n_4), .C(n_5), .Y(n_34) );
OAI222xp33_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_30), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_6), .Y(n_35) );
AND4x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_9), .C(n_12), .D(n_10), .Y(n_36) );
AND3x4_ASAP7_75t_L g37 ( .A(n_36), .B(n_32), .C(n_18), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_18), .B1(n_36), .B2(n_35), .Y(n_38) );
endmodule