module fake_jpeg_25955_n_93 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_37),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_40),
.B1(n_38),
.B2(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_46),
.Y(n_60)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_65),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_48),
.B1(n_41),
.B2(n_39),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B(n_18),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_0),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_43),
.C(n_51),
.Y(n_65)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_74),
.B1(n_64),
.B2(n_66),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_20),
.A3(n_36),
.B1(n_35),
.B2(n_5),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_67),
.B1(n_2),
.B2(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_69),
.B1(n_3),
.B2(n_2),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_6),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_77),
.B(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_78),
.B1(n_14),
.B2(n_15),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_16),
.B1(n_17),
.B2(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_28),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_29),
.C(n_30),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_31),
.B(n_32),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_33),
.Y(n_93)
);


endmodule