module fake_jpeg_25231_n_33 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx13_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_3),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_10),
.B1(n_8),
.B2(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_15),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_10),
.C(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_19),
.Y(n_23)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_20),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_23),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_25),
.C(n_18),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_28),
.A3(n_22),
.B1(n_11),
.B2(n_18),
.C1(n_15),
.C2(n_14),
.Y(n_31)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_11),
.CI(n_5),
.CON(n_32),
.SN(n_32)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_1),
.B(n_9),
.Y(n_33)
);


endmodule