module real_jpeg_25365_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_286;
wire n_176;
wire n_292;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_216;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_2),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_22),
.B1(n_51),
.B2(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_22),
.B1(n_71),
.B2(n_72),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_19),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_5),
.A2(n_32),
.B1(n_51),
.B2(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_32),
.B1(n_71),
.B2(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_58),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_20),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_41),
.B1(n_71),
.B2(n_72),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_26),
.C(n_30),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_8),
.B(n_27),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_8),
.B(n_48),
.C(n_51),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_8),
.B(n_68),
.C(n_71),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_8),
.B(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_8),
.B(n_102),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_8),
.B(n_61),
.Y(n_251)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_74),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_34),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_34),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_17),
.A2(n_37),
.B(n_38),
.Y(n_36)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_19),
.B(n_188),
.Y(n_187)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_23),
.A2(n_27),
.B1(n_39),
.B2(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_30),
.B(n_223),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_35),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_35),
.B(n_291),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_42),
.CI(n_54),
.CON(n_35),
.SN(n_35)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_37),
.A2(n_38),
.B(n_57),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_45),
.A2(n_50),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_61),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_46),
.B(n_107),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_50),
.A2(n_106),
.B(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_51),
.B(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_62),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_55),
.B(n_125),
.C(n_133),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_55),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_55),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_133),
.B1(n_134),
.B2(n_147),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_55),
.A2(n_104),
.B1(n_147),
.B2(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_55),
.B(n_104),
.C(n_185),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_59),
.A2(n_62),
.B1(n_114),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_59),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_62),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_62),
.B(n_110),
.C(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_73),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_64),
.B(n_92),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_66),
.A2(n_92),
.B1(n_102),
.B2(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_70),
.A2(n_91),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_71),
.B(n_241),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_290),
.B(n_292),
.Y(n_76)
);

OAI211xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_135),
.B(n_149),
.C(n_289),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_119),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_119),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_97),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_99),
.C(n_108),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_88),
.B(n_93),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_93),
.B1(n_94),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_89),
.B1(n_122),
.B2(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_83),
.B(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_87),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_86),
.A2(n_127),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_86),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_89),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_108),
.B2(n_109),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_100),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_207),
.C(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_104),
.A2(n_197),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_111),
.B1(n_143),
.B2(n_148),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_133),
.C(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_110),
.A2(n_111),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_110),
.A2(n_111),
.B1(n_167),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_159),
.C(n_167),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_111),
.B(n_139),
.C(n_143),
.Y(n_291)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_123),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_126),
.Y(n_280)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_130),
.A2(n_131),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_130),
.A2(n_131),
.B1(n_220),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_214),
.C(n_220),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_131),
.B(n_190),
.C(n_251),
.Y(n_255)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_133),
.A2(n_134),
.B1(n_181),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_133),
.A2(n_134),
.B1(n_165),
.B2(n_178),
.Y(n_257)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_134),
.B(n_165),
.C(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_150),
.C(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_137),
.B(n_138),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_171),
.B(n_288),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_169),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_153),
.B(n_169),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_158),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_154),
.B(n_156),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_158),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_159),
.A2(n_160),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_165),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_192),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_165),
.A2(n_178),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_283),
.B(n_287),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_210),
.B(n_269),
.C(n_282),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_199),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_199),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_184),
.B2(n_198),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_177),
.B(n_183),
.C(n_198),
.Y(n_270)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_189),
.A2(n_190),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_243),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_190)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_201),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_208),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_268),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_229),
.B(n_267),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_226),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_226),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_215),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_260),
.B(n_266),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_254),
.B(n_259),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_246),
.B(n_253),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_245),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_242),
.B(n_244),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_278),
.B2(n_279),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_279),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);


endmodule