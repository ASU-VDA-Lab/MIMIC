module fake_jpeg_26169_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_45),
.B1(n_16),
.B2(n_25),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_46),
.B(n_33),
.C(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_34),
.C(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_25),
.B1(n_19),
.B2(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_32),
.B1(n_22),
.B2(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_16),
.B1(n_13),
.B2(n_18),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22x1_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_30),
.B1(n_15),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_32),
.B(n_30),
.C(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_20),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_44),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_32),
.B1(n_44),
.B2(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_18),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_30),
.B(n_31),
.C(n_29),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_35),
.A3(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_74),
.B1(n_52),
.B2(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_15),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_43),
.B1(n_64),
.B2(n_73),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.C(n_0),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_51),
.C(n_59),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_83),
.B(n_88),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_61),
.B(n_26),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_15),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_12),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_73),
.A3(n_29),
.B1(n_19),
.B2(n_40),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_97),
.B(n_83),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_43),
.B1(n_27),
.B2(n_47),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_19),
.B1(n_36),
.B2(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_36),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_76),
.C(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_81),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_93),
.B1(n_97),
.B2(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_77),
.C(n_9),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_11),
.C(n_10),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_91),
.A3(n_97),
.B1(n_90),
.B2(n_94),
.C1(n_98),
.C2(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_110),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_103),
.B(n_102),
.Y(n_122)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_109),
.B(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_118),
.C(n_10),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_9),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_118),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_130),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_128),
.B1(n_125),
.B2(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_3),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_124),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_6),
.B(n_133),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_134),
.B(n_5),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_5),
.B(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_6),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_138),
.CI(n_129),
.CON(n_141),
.SN(n_141)
);


endmodule