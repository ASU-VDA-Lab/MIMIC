module fake_jpeg_13090_n_514 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_51),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_71),
.Y(n_133)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_69),
.Y(n_122)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_8),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_92),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_17),
.B1(n_7),
.B2(n_9),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_34),
.B1(n_31),
.B2(n_42),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_38),
.B(n_6),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_107),
.B(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_26),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_53),
.B1(n_58),
.B2(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_117),
.A2(n_157),
.B1(n_50),
.B2(n_97),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_119),
.A2(n_161),
.B1(n_6),
.B2(n_15),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_32),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_63),
.A2(n_49),
.B1(n_37),
.B2(n_45),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_123),
.A2(n_125),
.B(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_55),
.A2(n_37),
.B1(n_18),
.B2(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_60),
.A2(n_18),
.B1(n_37),
.B2(n_43),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_126),
.A2(n_66),
.B1(n_28),
.B2(n_91),
.Y(n_195)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_55),
.A2(n_18),
.B1(n_43),
.B2(n_28),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_59),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_67),
.A2(n_42),
.B1(n_30),
.B2(n_31),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_72),
.A2(n_30),
.B1(n_44),
.B2(n_36),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_185),
.Y(n_222)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_50),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_203),
.Y(n_257)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_79),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_174),
.B(n_183),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_184),
.C(n_207),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_36),
.B1(n_44),
.B2(n_78),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_101),
.B(n_116),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_189),
.C(n_205),
.Y(n_227)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_79),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_103),
.B(n_138),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_135),
.B(n_130),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_196),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_66),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_114),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g272 ( 
.A(n_193),
.B(n_13),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_198),
.B1(n_162),
.B2(n_150),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_197),
.A2(n_5),
.B1(n_13),
.B2(n_12),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_125),
.A2(n_87),
.B1(n_75),
.B2(n_73),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_117),
.A2(n_152),
.B1(n_147),
.B2(n_134),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_200),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_0),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_156),
.B(n_28),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_120),
.A2(n_28),
.B1(n_51),
.B2(n_93),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_0),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_221),
.C(n_148),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_216),
.Y(n_243)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_218),
.Y(n_249)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_5),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_139),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_162),
.B1(n_134),
.B2(n_140),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_132),
.B(n_0),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_143),
.B(n_108),
.C(n_132),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_224),
.A2(n_185),
.B(n_209),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_248),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_234),
.A2(n_253),
.B1(n_270),
.B2(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_242),
.A2(n_268),
.B1(n_271),
.B2(n_273),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_170),
.A2(n_11),
.B(n_17),
.C(n_15),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_177),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_250),
.B(n_179),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_199),
.A2(n_155),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_258),
.B1(n_260),
.B2(n_168),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_179),
.B(n_3),
.C(n_4),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_221),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_214),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_202),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_167),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_165),
.B(n_17),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_269),
.B(n_173),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_210),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_272),
.A2(n_263),
.B(n_246),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_211),
.A2(n_212),
.B1(n_206),
.B2(n_193),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_274),
.A2(n_278),
.B1(n_285),
.B2(n_256),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_214),
.B(n_221),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_277),
.A2(n_291),
.B(n_310),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_234),
.A2(n_219),
.B1(n_205),
.B2(n_203),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_279),
.B(n_237),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_284),
.C(n_299),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_303),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_257),
.B(n_182),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_282),
.B(n_304),
.Y(n_328)
);

BUFx4f_ASAP7_75t_SL g283 ( 
.A(n_231),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_181),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_204),
.B1(n_218),
.B2(n_191),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_259),
.A2(n_216),
.B1(n_194),
.B2(n_208),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_171),
.B(n_172),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_294),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_180),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_302),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_297),
.B1(n_315),
.B2(n_266),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_190),
.B1(n_169),
.B2(n_163),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_227),
.B(n_178),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_225),
.Y(n_300)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_222),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_192),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_305),
.B(n_312),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_259),
.A2(n_166),
.B1(n_217),
.B2(n_245),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_309),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_240),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_318),
.Y(n_355)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_241),
.B(n_227),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_224),
.A2(n_272),
.B(n_270),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_313),
.B(n_246),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_241),
.B(n_230),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_235),
.B(n_233),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_316),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_260),
.B1(n_253),
.B2(n_233),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_266),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_320),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_265),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_296),
.A2(n_310),
.B1(n_315),
.B2(n_311),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_324),
.A2(n_325),
.B1(n_340),
.B2(n_346),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_291),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_338),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_267),
.B1(n_232),
.B2(n_265),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_237),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_280),
.C(n_298),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_314),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_310),
.A2(n_232),
.B1(n_267),
.B2(n_247),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_342),
.B(n_353),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_322),
.B(n_336),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_262),
.B1(n_244),
.B2(n_226),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_317),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_338),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_294),
.A2(n_262),
.B1(n_244),
.B2(n_226),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_357),
.B1(n_276),
.B2(n_293),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_281),
.A2(n_285),
.B1(n_308),
.B2(n_282),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_352),
.A2(n_356),
.B1(n_301),
.B2(n_304),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_284),
.B(n_256),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_295),
.A2(n_229),
.B1(n_239),
.B2(n_254),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_322),
.A2(n_305),
.B1(n_275),
.B2(n_286),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_362),
.A2(n_363),
.B(n_367),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_288),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_374),
.B(n_379),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_355),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_359),
.A2(n_277),
.B1(n_298),
.B2(n_289),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_370),
.C(n_371),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_369),
.A2(n_377),
.B1(n_329),
.B2(n_385),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_279),
.C(n_313),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

A2O1A1O1Ixp25_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_320),
.B(n_254),
.C(n_302),
.D(n_292),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_331),
.A2(n_309),
.B(n_307),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_363),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_343),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_290),
.B(n_251),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_391),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_319),
.B(n_318),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_356),
.A2(n_300),
.B1(n_239),
.B2(n_229),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_381),
.A2(n_382),
.B1(n_329),
.B2(n_378),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_333),
.A2(n_251),
.B1(n_283),
.B2(n_325),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_283),
.Y(n_383)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_283),
.C(n_342),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_386),
.C(n_393),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_333),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_360),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_337),
.A2(n_339),
.B(n_327),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_339),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_327),
.A2(n_360),
.B1(n_346),
.B2(n_326),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_349),
.B1(n_341),
.B2(n_348),
.Y(n_406)
);

AOI221xp5_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_354),
.B1(n_358),
.B2(n_330),
.C(n_349),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_396),
.B(n_374),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_330),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_380),
.Y(n_402)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_406),
.A2(n_410),
.B1(n_421),
.B2(n_407),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_361),
.A2(n_341),
.B1(n_343),
.B2(n_348),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_415),
.B1(n_421),
.B2(n_385),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_321),
.Y(n_409)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

AOI211xp5_ASAP7_75t_SL g410 ( 
.A1(n_363),
.A2(n_321),
.B(n_329),
.C(n_364),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_412),
.A2(n_414),
.B1(n_390),
.B2(n_379),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_361),
.A2(n_362),
.B1(n_373),
.B2(n_394),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_370),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_393),
.C(n_391),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_417),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_373),
.A2(n_366),
.B1(n_363),
.B2(n_367),
.Y(n_421)
);

FAx1_ASAP7_75t_SL g423 ( 
.A(n_368),
.B(n_388),
.CI(n_384),
.CON(n_423),
.SN(n_423)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_386),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_424),
.B(n_425),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_431),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_428),
.B(n_439),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_416),
.C(n_405),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_438),
.C(n_397),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_430),
.A2(n_441),
.B1(n_419),
.B2(n_420),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_376),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_402),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_444),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_390),
.B1(n_378),
.B2(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_443),
.B1(n_446),
.B2(n_417),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_381),
.Y(n_436)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_398),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_423),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_401),
.C(n_395),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_413),
.B(n_418),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_400),
.A2(n_413),
.B(n_403),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_433),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_395),
.A2(n_404),
.B1(n_400),
.B2(n_403),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_408),
.B(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_404),
.B1(n_408),
.B2(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_412),
.Y(n_447)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_447),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_399),
.B(n_397),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_462),
.B(n_455),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_442),
.B1(n_427),
.B2(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_456),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_463),
.B(n_448),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_458),
.A2(n_462),
.B1(n_454),
.B2(n_465),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_431),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_459),
.B(n_460),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_425),
.C(n_426),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_433),
.B(n_435),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_441),
.Y(n_463)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_463),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_447),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_455),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_442),
.Y(n_469)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_437),
.C(n_424),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_472),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_460),
.C(n_456),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_449),
.Y(n_474)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_476),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_SL g483 ( 
.A(n_477),
.B(n_479),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_450),
.C(n_458),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_481),
.B(n_461),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_457),
.C(n_464),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_472),
.C(n_480),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_487),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_452),
.C(n_449),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_490),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_475),
.A2(n_469),
.B(n_468),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_476),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_482),
.B(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_495),
.Y(n_501)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_485),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_477),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_491),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_492),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_500),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_484),
.A2(n_486),
.B1(n_473),
.B2(n_470),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_491),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_493),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_496),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_499),
.B(n_498),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_507),
.B(n_483),
.Y(n_509)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_506),
.A2(n_504),
.B(n_474),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_508),
.A2(n_509),
.B(n_494),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_510),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_489),
.B(n_502),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_478),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_513),
.B(n_471),
.Y(n_514)
);


endmodule