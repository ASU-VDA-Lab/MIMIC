module real_aes_4155_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_617;
wire n_733;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_483;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_0), .A2(n_287), .B1(n_561), .B2(n_570), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_1), .A2(n_401), .B1(n_564), .B2(n_565), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_2), .A2(n_6), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_3), .A2(n_91), .B1(n_530), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_4), .A2(n_69), .B1(n_729), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_5), .A2(n_216), .B1(n_562), .B2(n_568), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_7), .A2(n_179), .B1(n_723), .B2(n_728), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_8), .A2(n_360), .B1(n_562), .B2(n_568), .Y(n_746) );
INVx1_ASAP7_75t_L g781 ( .A(n_9), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_10), .A2(n_309), .B1(n_1062), .B2(n_1342), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_11), .A2(n_106), .B1(n_671), .B2(n_729), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_12), .A2(n_183), .B1(n_651), .B2(n_801), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_13), .A2(n_52), .B1(n_679), .B2(n_726), .Y(n_765) );
AOI21x1_ASAP7_75t_L g775 ( .A1(n_14), .A2(n_776), .B(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g840 ( .A(n_15), .Y(n_840) );
INVx1_ASAP7_75t_SL g1201 ( .A(n_16), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_17), .A2(n_379), .B1(n_723), .B2(n_865), .Y(n_1038) );
INVx1_ASAP7_75t_L g859 ( .A(n_18), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_19), .A2(n_341), .B1(n_446), .B2(n_490), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_20), .A2(n_36), .B1(n_677), .B2(n_767), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_21), .A2(n_109), .B1(n_723), .B2(n_883), .Y(n_1008) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_22), .B(n_452), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_23), .A2(n_290), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g1108 ( .A(n_24), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_25), .A2(n_270), .B1(n_564), .B2(n_565), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_26), .A2(n_186), .B1(n_627), .B2(n_883), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_27), .B(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_28), .A2(n_227), .B1(n_548), .B2(n_571), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_29), .A2(n_260), .B1(n_530), .B2(n_532), .Y(n_867) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_30), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_31), .A2(n_113), .B1(n_1095), .B2(n_1117), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_32), .A2(n_82), .B1(n_814), .B2(n_816), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_33), .A2(n_165), .B1(n_729), .B2(n_762), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_34), .A2(n_890), .B(n_891), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_35), .A2(n_48), .B1(n_670), .B2(n_672), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_37), .A2(n_157), .B1(n_538), .B2(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g797 ( .A(n_38), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_39), .A2(n_234), .B1(n_549), .B2(n_554), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_40), .A2(n_304), .B1(n_864), .B2(n_865), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_41), .B(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_42), .A2(n_261), .B1(n_1135), .B2(n_1138), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_43), .A2(n_114), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g1360 ( .A1(n_44), .A2(n_1361), .B1(n_1362), .B2(n_1378), .Y(n_1360) );
INVx1_ASAP7_75t_L g1378 ( .A(n_44), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_45), .A2(n_226), .B1(n_676), .B2(n_677), .Y(n_978) );
XOR2x2_ASAP7_75t_L g987 ( .A(n_46), .B(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_47), .A2(n_405), .B1(n_549), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_49), .A2(n_163), .B1(n_532), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1104 ( .A(n_50), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_51), .A2(n_121), .B1(n_486), .B2(n_490), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_53), .A2(n_145), .B1(n_486), .B2(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g905 ( .A(n_54), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_55), .A2(n_354), .B1(n_624), .B2(n_627), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_56), .A2(n_104), .B1(n_511), .B2(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g637 ( .A(n_57), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_58), .A2(n_154), .B1(n_530), .B2(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_59), .A2(n_180), .B1(n_647), .B2(n_671), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_60), .A2(n_200), .B1(n_536), .B2(n_655), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_61), .B(n_704), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_62), .A2(n_118), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_63), .A2(n_257), .B1(n_562), .B2(n_568), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_64), .A2(n_282), .B1(n_567), .B2(n_582), .Y(n_581) );
OA22x2_ASAP7_75t_L g467 ( .A1(n_65), .A2(n_177), .B1(n_452), .B2(n_466), .Y(n_467) );
INVx1_ASAP7_75t_L g496 ( .A(n_65), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_66), .A2(n_348), .B1(n_673), .B2(n_762), .Y(n_898) );
XNOR2x1_ASAP7_75t_L g874 ( .A(n_67), .B(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_68), .A2(n_75), .B1(n_703), .B2(n_704), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_70), .A2(n_72), .B1(n_564), .B2(n_565), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_71), .A2(n_334), .B1(n_526), .B2(n_864), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_73), .A2(n_400), .B1(n_663), .B2(n_857), .Y(n_1045) );
XNOR2x2_ASAP7_75t_L g919 ( .A(n_74), .B(n_920), .Y(n_919) );
XOR2x2_ASAP7_75t_L g758 ( .A(n_76), .B(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_77), .A2(n_278), .B1(n_551), .B2(n_552), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_78), .A2(n_340), .B1(n_564), .B2(n_565), .Y(n_1033) );
INVx1_ASAP7_75t_L g715 ( .A(n_79), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_80), .A2(n_117), .B1(n_522), .B2(n_526), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_81), .A2(n_289), .B1(n_548), .B2(n_571), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_83), .A2(n_208), .B1(n_819), .B2(n_845), .C(n_990), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_84), .B(n_202), .Y(n_432) );
INVx1_ASAP7_75t_L g465 ( .A(n_84), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_84), .A2(n_177), .B(n_478), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g810 ( .A1(n_85), .A2(n_499), .B(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_86), .A2(n_166), .B1(n_714), .B2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_87), .A2(n_396), .B1(n_564), .B2(n_565), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_88), .A2(n_134), .B1(n_767), .B2(n_768), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_89), .A2(n_306), .B1(n_624), .B2(n_627), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_90), .A2(n_159), .B1(n_511), .B2(n_729), .Y(n_973) );
INVx1_ASAP7_75t_L g1029 ( .A(n_92), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_93), .A2(n_194), .B1(n_1074), .B2(n_1352), .Y(n_1351) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_94), .A2(n_206), .B1(n_511), .B2(n_518), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_95), .A2(n_238), .B1(n_511), .B2(n_729), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_96), .A2(n_167), .B1(n_582), .B2(n_821), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_97), .A2(n_137), .B1(n_676), .B2(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_98), .B(n_861), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_99), .B(n_663), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_100), .A2(n_389), .B1(n_694), .B2(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g1097 ( .A(n_101), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_101), .B(n_302), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_102), .A2(n_355), .B1(n_548), .B2(n_571), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_103), .A2(n_263), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_105), .A2(n_224), .B1(n_582), .B2(n_741), .Y(n_1370) );
INVx1_ASAP7_75t_L g1051 ( .A(n_107), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_108), .A2(n_243), .B1(n_723), .B2(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_110), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_111), .A2(n_112), .B1(n_726), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g1081 ( .A(n_115), .Y(n_1081) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_116), .A2(n_120), .B1(n_694), .B2(n_1047), .C(n_1049), .Y(n_1046) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_119), .A2(n_567), .B(n_904), .Y(n_903) );
XNOR2x1_ASAP7_75t_L g709 ( .A(n_122), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_123), .A2(n_361), .B1(n_567), .B2(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_124), .B(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_125), .A2(n_170), .B1(n_536), .B2(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_126), .A2(n_222), .B1(n_486), .B2(n_490), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_127), .A2(n_171), .B1(n_530), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_128), .A2(n_201), .B1(n_549), .B2(n_552), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1374 ( .A1(n_129), .A2(n_160), .B1(n_1342), .B2(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1050 ( .A(n_130), .Y(n_1050) );
INVx1_ASAP7_75t_SL g1098 ( .A(n_131), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_131), .B(n_428), .Y(n_1101) );
INVx1_ASAP7_75t_L g1112 ( .A(n_131), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_132), .A2(n_286), .B1(n_490), .B2(n_597), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_133), .A2(n_193), .B1(n_645), .B2(n_648), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_135), .A2(n_213), .B1(n_751), .B2(n_928), .Y(n_927) );
XNOR2x1_ASAP7_75t_L g824 ( .A(n_136), .B(n_825), .Y(n_824) );
XNOR2x2_ASAP7_75t_SL g912 ( .A(n_136), .B(n_825), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_138), .A2(n_312), .B1(n_624), .B2(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g749 ( .A(n_139), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g1132 ( .A(n_140), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_141), .A2(n_168), .B1(n_1125), .B2(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g955 ( .A(n_142), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_143), .A2(n_292), .B1(n_530), .B2(n_532), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_144), .A2(n_399), .B1(n_551), .B2(n_567), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_146), .A2(n_409), .B1(n_844), .B2(n_845), .C(n_846), .Y(n_843) );
INVx1_ASAP7_75t_L g1099 ( .A(n_147), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_148), .A2(n_383), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_149), .A2(n_318), .B1(n_490), .B2(n_611), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_150), .A2(n_164), .B1(n_526), .B2(n_723), .Y(n_933) );
INVx1_ASAP7_75t_L g1348 ( .A(n_151), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_152), .A2(n_220), .B1(n_499), .B2(n_714), .Y(n_1014) );
OAI22x1_ASAP7_75t_L g961 ( .A1(n_153), .A2(n_962), .B1(n_984), .B2(n_985), .Y(n_961) );
NAND3xp33_ASAP7_75t_SL g984 ( .A(n_153), .B(n_972), .C(n_979), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_155), .A2(n_198), .B1(n_561), .B2(n_570), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_156), .A2(n_406), .B1(n_564), .B2(n_565), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_158), .A2(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g835 ( .A(n_161), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_162), .A2(n_190), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_169), .A2(n_251), .B1(n_1068), .B2(n_1334), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_172), .A2(n_244), .B1(n_714), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_173), .A2(n_339), .B1(n_538), .B2(n_880), .Y(n_942) );
CKINVDCx6p67_ASAP7_75t_R g1131 ( .A(n_174), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_175), .A2(n_392), .B1(n_548), .B2(n_571), .Y(n_744) );
INVx1_ASAP7_75t_L g459 ( .A(n_176), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_176), .B(n_242), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_176), .B(n_494), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_177), .B(n_317), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_178), .A2(n_252), .B1(n_536), .B2(n_538), .Y(n_866) );
INVx1_ASAP7_75t_L g812 ( .A(n_181), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_182), .A2(n_310), .B1(n_446), .B2(n_855), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_184), .A2(n_285), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_185), .A2(n_203), .B1(n_694), .B2(n_731), .C(n_733), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_187), .A2(n_347), .B1(n_536), .B2(n_538), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_188), .A2(n_195), .B1(n_446), .B2(n_783), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_189), .A2(n_265), .B1(n_536), .B2(n_538), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_191), .A2(n_352), .B1(n_670), .B2(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g502 ( .A(n_192), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_196), .A2(n_374), .B1(n_1106), .B2(n_1110), .Y(n_1118) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_197), .A2(n_546), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_199), .B(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_202), .B(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_204), .A2(n_235), .B1(n_532), .B2(n_647), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_205), .A2(n_284), .B1(n_561), .B2(n_570), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_207), .A2(n_419), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_209), .A2(n_250), .B1(n_671), .B2(n_729), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_210), .A2(n_420), .B1(n_538), .B2(n_726), .Y(n_725) );
AO22x2_ASAP7_75t_L g593 ( .A1(n_211), .A2(n_594), .B1(n_617), .B2(n_618), .Y(n_593) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_211), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_211), .A2(n_323), .B1(n_1106), .B2(n_1110), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_212), .A2(n_273), .B1(n_814), .B2(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g892 ( .A(n_214), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_215), .A2(n_338), .B1(n_530), .B2(n_936), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_217), .B(n_606), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_218), .B(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_219), .A2(n_394), .B1(n_446), .B2(n_468), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_221), .A2(n_939), .B1(n_940), .B2(n_956), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_221), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_223), .A2(n_344), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_225), .A2(n_255), .B1(n_694), .B2(n_816), .Y(n_1015) );
XNOR2x1_ASAP7_75t_L g895 ( .A(n_228), .B(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_229), .A2(n_417), .B1(n_538), .B2(n_880), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_230), .A2(n_410), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
BUFx2_ASAP7_75t_L g604 ( .A(n_231), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_232), .A2(n_275), .B1(n_864), .B2(n_1337), .Y(n_1336) );
XNOR2x1_ASAP7_75t_L g850 ( .A(n_233), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g632 ( .A(n_236), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g1116 ( .A1(n_237), .A2(n_391), .B1(n_1095), .B2(n_1117), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_239), .A2(n_313), .B1(n_1122), .B2(n_1138), .Y(n_1161) );
INVx1_ASAP7_75t_L g734 ( .A(n_240), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_241), .A2(n_421), .B1(n_499), .B2(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g463 ( .A(n_242), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_245), .B(n_966), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_246), .A2(n_416), .B1(n_651), .B2(n_679), .Y(n_678) );
XNOR2x1_ASAP7_75t_L g542 ( .A(n_247), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_247), .A2(n_259), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_248), .A2(n_386), .B1(n_821), .B2(n_822), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_249), .A2(n_384), .B1(n_446), .B2(n_857), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_253), .A2(n_264), .B1(n_714), .B2(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_254), .B(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_256), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_258), .A2(n_366), .B1(n_522), .B2(n_865), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_262), .A2(n_331), .B1(n_627), .B2(n_936), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_266), .A2(n_320), .B1(n_647), .B2(n_947), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_267), .A2(n_288), .B1(n_561), .B2(n_570), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_268), .A2(n_350), .B1(n_511), .B2(n_829), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_269), .A2(n_330), .B1(n_562), .B2(n_568), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_271), .A2(n_298), .B1(n_1125), .B2(n_1126), .Y(n_1147) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_272), .B(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_274), .A2(n_356), .B1(n_499), .B2(n_1368), .Y(n_1367) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_276), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_277), .A2(n_325), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_279), .A2(n_315), .B1(n_783), .B2(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_280), .A2(n_326), .B1(n_532), .B2(n_647), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_281), .A2(n_357), .B1(n_651), .B2(n_654), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_283), .A2(n_398), .B1(n_649), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_291), .A2(n_308), .B1(n_551), .B2(n_552), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_293), .A2(n_415), .B1(n_1352), .B2(n_1366), .Y(n_1365) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_294), .A2(n_296), .B1(n_741), .B2(n_1077), .C(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g784 ( .A(n_295), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_297), .A2(n_342), .B1(n_561), .B2(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g842 ( .A(n_299), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_300), .A2(n_324), .B1(n_1123), .B2(n_1135), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1353 ( .A1(n_301), .A2(n_335), .B1(n_980), .B2(n_1071), .Y(n_1353) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_302), .Y(n_433) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_302), .B(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_303), .B(n_731), .Y(n_952) );
XNOR2x2_ASAP7_75t_L g1055 ( .A(n_305), .B(n_1056), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_307), .A2(n_346), .B1(n_561), .B2(n_570), .Y(n_1034) );
INVx1_ASAP7_75t_L g716 ( .A(n_311), .Y(n_716) );
XOR2x2_ASAP7_75t_L g620 ( .A(n_313), .B(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_314), .A2(n_371), .B1(n_549), .B2(n_567), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_316), .A2(n_337), .B1(n_627), .B2(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g457 ( .A(n_317), .Y(n_457) );
INVxp67_ASAP7_75t_L g477 ( .A(n_317), .Y(n_477) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_319), .A2(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g991 ( .A(n_321), .Y(n_991) );
INVx1_ASAP7_75t_L g755 ( .A(n_322), .Y(n_755) );
INVx1_ASAP7_75t_L g573 ( .A(n_324), .Y(n_573) );
AOI22xp5_ASAP7_75t_SL g979 ( .A1(n_327), .A2(n_381), .B1(n_980), .B2(n_982), .Y(n_979) );
INVxp67_ASAP7_75t_R g1136 ( .A(n_328), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_329), .A2(n_349), .B1(n_562), .B2(n_568), .Y(n_1032) );
INVx2_ASAP7_75t_L g428 ( .A(n_332), .Y(n_428) );
INVx1_ASAP7_75t_L g634 ( .A(n_333), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_336), .A2(n_923), .B(n_924), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_343), .A2(n_345), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g658 ( .A(n_351), .Y(n_658) );
INVx1_ASAP7_75t_L g639 ( .A(n_353), .Y(n_639) );
INVx1_ASAP7_75t_L g847 ( .A(n_358), .Y(n_847) );
INVx1_ASAP7_75t_L g599 ( .A(n_359), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_362), .A2(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_363), .Y(n_556) );
INVx1_ASAP7_75t_L g718 ( .A(n_364), .Y(n_718) );
AOI21xp33_ASAP7_75t_SL g1344 ( .A1(n_365), .A2(n_1345), .B(n_1347), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_367), .B(n_660), .Y(n_1369) );
AOI21xp33_ASAP7_75t_L g856 ( .A1(n_368), .A2(n_857), .B(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_369), .A2(n_373), .B1(n_649), .B2(n_673), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_370), .A2(n_408), .B1(n_651), .B2(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_372), .A2(n_390), .B1(n_490), .B2(n_611), .Y(n_906) );
INVx1_ASAP7_75t_L g442 ( .A(n_374), .Y(n_442) );
INVx1_ASAP7_75t_L g1102 ( .A(n_375), .Y(n_1102) );
OAI22x1_ASAP7_75t_L g1329 ( .A1(n_375), .A2(n_1102), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_375), .A2(n_1359), .B1(n_1379), .B2(n_1381), .Y(n_1358) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_376), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_377), .A2(n_413), .B1(n_548), .B2(n_571), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_378), .B(n_664), .Y(n_926) );
INVx1_ASAP7_75t_L g1021 ( .A(n_380), .Y(n_1021) );
XNOR2x2_ASAP7_75t_L g667 ( .A(n_382), .B(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_385), .A2(n_404), .B1(n_624), .B2(n_627), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_387), .A2(n_412), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
INVx1_ASAP7_75t_SL g1018 ( .A(n_388), .Y(n_1018) );
INVx1_ASAP7_75t_L g756 ( .A(n_393), .Y(n_756) );
BUFx2_ASAP7_75t_L g608 ( .A(n_395), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_397), .B(n_579), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_402), .A2(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g1202 ( .A(n_403), .Y(n_1202) );
INVx1_ASAP7_75t_L g925 ( .A(n_407), .Y(n_925) );
AOI21xp33_ASAP7_75t_L g1027 ( .A1(n_411), .A2(n_554), .B(n_1028), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_414), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g953 ( .A1(n_418), .A2(n_930), .B(n_954), .Y(n_953) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_434), .B(n_1083), .Y(n_422) );
INVx2_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
BUFx4_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .C(n_433), .Y(n_425) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_426), .B(n_1356), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_426), .B(n_1357), .Y(n_1380) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OA21x2_ASAP7_75t_L g1382 ( .A1(n_427), .A2(n_1098), .B(n_1383), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND3x4_ASAP7_75t_L g1095 ( .A(n_428), .B(n_1096), .C(n_1098), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_428), .B(n_1112), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_429), .B(n_1357), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_430), .A2(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g1357 ( .A(n_433), .Y(n_1357) );
XNOR2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_790), .Y(n_434) );
XNOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_666), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_589), .B2(n_665), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
XOR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_540), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
XOR2xp5_ASAP7_75t_L g592 ( .A(n_441), .B(n_593), .Y(n_592) );
XNOR2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_444), .B(n_509), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_479), .C(n_485), .D(n_498), .Y(n_444) );
INVx2_ASAP7_75t_L g981 ( .A(n_446), .Y(n_981) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_446), .Y(n_1072) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g642 ( .A(n_447), .Y(n_642) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_447), .Y(n_714) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
AND2x4_ASAP7_75t_L g500 ( .A(n_448), .B(n_488), .Y(n_500) );
AND2x4_ASAP7_75t_L g537 ( .A(n_448), .B(n_513), .Y(n_537) );
AND2x4_ASAP7_75t_L g551 ( .A(n_448), .B(n_460), .Y(n_551) );
AND2x4_ASAP7_75t_L g564 ( .A(n_448), .B(n_513), .Y(n_564) );
AND2x4_ASAP7_75t_L g567 ( .A(n_448), .B(n_488), .Y(n_567) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_454), .Y(n_448) );
AND2x2_ASAP7_75t_L g471 ( .A(n_449), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g484 ( .A(n_449), .Y(n_484) );
OR2x2_ASAP7_75t_L g516 ( .A(n_449), .B(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g524 ( .A(n_449), .B(n_525), .Y(n_524) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_451), .B(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g494 ( .A(n_451), .Y(n_494) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp33_ASAP7_75t_L g458 ( .A(n_452), .B(n_459), .Y(n_458) );
NAND2xp33_ASAP7_75t_L g462 ( .A(n_452), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_452), .Y(n_473) );
INVx1_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_453), .B(n_493), .C(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g483 ( .A(n_454), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
AND2x2_ASAP7_75t_L g482 ( .A(n_460), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g523 ( .A(n_460), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g527 ( .A(n_460), .B(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g562 ( .A(n_460), .B(n_515), .Y(n_562) );
AND2x4_ASAP7_75t_L g568 ( .A(n_460), .B(n_524), .Y(n_568) );
AND2x2_ASAP7_75t_L g628 ( .A(n_460), .B(n_524), .Y(n_628) );
AND2x2_ASAP7_75t_L g753 ( .A(n_460), .B(n_483), .Y(n_753) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_467), .Y(n_460) );
INVx1_ASAP7_75t_L g489 ( .A(n_461), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_463), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_465), .A2(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g475 ( .A(n_467), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g488 ( .A(n_467), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g514 ( .A(n_467), .Y(n_514) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g703 ( .A(n_469), .Y(n_703) );
INVx3_ASAP7_75t_L g741 ( .A(n_469), .Y(n_741) );
INVx4_ASAP7_75t_L g783 ( .A(n_469), .Y(n_783) );
INVx2_ASAP7_75t_L g821 ( .A(n_469), .Y(n_821) );
INVx5_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx4f_ASAP7_75t_L g663 ( .A(n_470), .Y(n_663) );
BUFx2_ASAP7_75t_L g855 ( .A(n_470), .Y(n_855) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
AND2x2_ASAP7_75t_L g552 ( .A(n_471), .B(n_475), .Y(n_552) );
AND2x4_ASAP7_75t_L g606 ( .A(n_471), .B(n_475), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g506 ( .A(n_473), .Y(n_506) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_SL g701 ( .A(n_481), .Y(n_701) );
INVx2_ASAP7_75t_L g819 ( .A(n_481), .Y(n_819) );
INVx2_ASAP7_75t_L g861 ( .A(n_481), .Y(n_861) );
INVx2_ASAP7_75t_L g1079 ( .A(n_481), .Y(n_1079) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
INVx2_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
AND2x4_ASAP7_75t_L g487 ( .A(n_483), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g491 ( .A(n_483), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g539 ( .A(n_483), .B(n_513), .Y(n_539) );
AND2x4_ASAP7_75t_L g549 ( .A(n_483), .B(n_492), .Y(n_549) );
AND2x2_ASAP7_75t_L g554 ( .A(n_483), .B(n_488), .Y(n_554) );
AND2x4_ASAP7_75t_L g565 ( .A(n_483), .B(n_513), .Y(n_565) );
BUFx3_ASAP7_75t_L g1074 ( .A(n_486), .Y(n_1074) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_487), .Y(n_611) );
BUFx3_ASAP7_75t_L g694 ( .A(n_487), .Y(n_694) );
BUFx8_ASAP7_75t_SL g751 ( .A(n_487), .Y(n_751) );
INVx2_ASAP7_75t_L g815 ( .A(n_487), .Y(n_815) );
AND2x4_ASAP7_75t_L g513 ( .A(n_489), .B(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g635 ( .A(n_490), .Y(n_635) );
BUFx3_ASAP7_75t_L g697 ( .A(n_490), .Y(n_697) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g774 ( .A(n_491), .Y(n_774) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_491), .Y(n_816) );
AND2x4_ASAP7_75t_L g520 ( .A(n_492), .B(n_515), .Y(n_520) );
AND2x4_ASAP7_75t_L g534 ( .A(n_492), .B(n_524), .Y(n_534) );
AND2x4_ASAP7_75t_L g570 ( .A(n_492), .B(n_524), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_492), .B(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx4_ASAP7_75t_L g638 ( .A(n_499), .Y(n_638) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g597 ( .A(n_500), .Y(n_597) );
INVx1_ASAP7_75t_L g686 ( .A(n_500), .Y(n_686) );
BUFx3_ASAP7_75t_L g857 ( .A(n_500), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g786 ( .A(n_504), .Y(n_786) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_504), .Y(n_848) );
INVx1_ASAP7_75t_L g1017 ( .A(n_504), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
NAND4xp25_ASAP7_75t_SL g509 ( .A(n_510), .B(n_521), .C(n_529), .D(n_535), .Y(n_509) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_512), .Y(n_649) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_512), .Y(n_671) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_512), .Y(n_762) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
AND2x4_ASAP7_75t_L g531 ( .A(n_513), .B(n_524), .Y(n_531) );
AND2x4_ASAP7_75t_L g548 ( .A(n_513), .B(n_528), .Y(n_548) );
AND2x4_ASAP7_75t_L g561 ( .A(n_513), .B(n_524), .Y(n_561) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g528 ( .A(n_516), .Y(n_528) );
INVx1_ASAP7_75t_L g525 ( .A(n_517), .Y(n_525) );
BUFx2_ASAP7_75t_L g625 ( .A(n_518), .Y(n_625) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g673 ( .A(n_519), .Y(n_673) );
INVx3_ASAP7_75t_L g829 ( .A(n_519), .Y(n_829) );
INVx1_ASAP7_75t_L g878 ( .A(n_519), .Y(n_878) );
INVx1_ASAP7_75t_L g1373 ( .A(n_519), .Y(n_1373) );
INVx6_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx12f_ASAP7_75t_L g729 ( .A(n_520), .Y(n_729) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_523), .Y(n_864) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g624 ( .A(n_527), .Y(n_624) );
BUFx12f_ASAP7_75t_L g728 ( .A(n_527), .Y(n_728) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_527), .Y(n_865) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_527), .Y(n_883) );
BUFx2_ASAP7_75t_SL g1061 ( .A(n_530), .Y(n_1061) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx12f_ASAP7_75t_L g647 ( .A(n_531), .Y(n_647) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_531), .Y(n_767) );
BUFx2_ASAP7_75t_SL g1062 ( .A(n_532), .Y(n_1062) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g629 ( .A(n_533), .Y(n_629) );
INVx4_ASAP7_75t_L g677 ( .A(n_533), .Y(n_677) );
INVx1_ASAP7_75t_L g768 ( .A(n_533), .Y(n_768) );
INVx4_ASAP7_75t_L g885 ( .A(n_533), .Y(n_885) );
INVx4_ASAP7_75t_L g936 ( .A(n_533), .Y(n_936) );
INVx2_ASAP7_75t_L g947 ( .A(n_533), .Y(n_947) );
INVx8_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx12f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g653 ( .A(n_537), .Y(n_653) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_537), .Y(n_726) );
BUFx2_ASAP7_75t_SL g1340 ( .A(n_538), .Y(n_1340) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
BUFx5_ASAP7_75t_L g679 ( .A(n_539), .Y(n_679) );
INVx1_ASAP7_75t_L g803 ( .A(n_539), .Y(n_803) );
OA22x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_572), .B2(n_588), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
XOR2x2_ASAP7_75t_L g937 ( .A(n_542), .B(n_938), .Y(n_937) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_559), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .C(n_550), .D(n_553), .Y(n_544) );
INVx1_ASAP7_75t_L g661 ( .A(n_546), .Y(n_661) );
INVx2_ASAP7_75t_L g779 ( .A(n_546), .Y(n_779) );
BUFx3_ASAP7_75t_L g1346 ( .A(n_546), .Y(n_1346) );
INVx2_ASAP7_75t_L g841 ( .A(n_549), .Y(n_841) );
INVx2_ASAP7_75t_L g609 ( .A(n_551), .Y(n_609) );
INVx1_ASAP7_75t_L g839 ( .A(n_551), .Y(n_839) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_554), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g582 ( .A(n_557), .Y(n_582) );
INVx4_ASAP7_75t_L g664 ( .A(n_557), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_557), .B(n_991), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_557), .B(n_1029), .Y(n_1028) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g600 ( .A(n_558), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .C(n_566), .D(n_569), .Y(n_559) );
INVx2_ASAP7_75t_L g836 ( .A(n_567), .Y(n_836) );
XNOR2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
XOR2xp5_ASAP7_75t_L g588 ( .A(n_573), .B(n_574), .Y(n_588) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_583), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .C(n_578), .D(n_581), .Y(n_575) );
INVx1_ASAP7_75t_L g967 ( .A(n_579), .Y(n_967) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_580), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .C(n_586), .D(n_587), .Y(n_583) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g665 ( .A(n_590), .Y(n_665) );
AO22x2_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_619), .B2(n_620), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g618 ( .A(n_594), .Y(n_618) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_612), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_601), .C(n_610), .Y(n_595) );
INVx2_ASAP7_75t_L g983 ( .A(n_597), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx4_ASAP7_75t_L g704 ( .A(n_600), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_600), .B(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_600), .B(n_812), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_600), .B(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_600), .B(n_1050), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1080 ( .A(n_600), .B(n_1081), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B1(n_607), .B2(n_609), .Y(n_602) );
CKINVDCx16_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g891 ( .A1(n_605), .A2(n_892), .B(n_893), .Y(n_891) );
OAI21xp33_ASAP7_75t_L g924 ( .A1(n_605), .A2(n_925), .B(n_926), .Y(n_924) );
INVx4_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx9p33_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g633 ( .A(n_611), .Y(n_633) );
BUFx3_ASAP7_75t_L g1366 ( .A(n_611), .Y(n_1366) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .C(n_615), .D(n_616), .Y(n_612) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_630), .C(n_643), .D(n_656), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
BUFx8_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_628), .Y(n_723) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_636), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_635), .A2(n_713), .B1(n_715), .B2(n_716), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_638), .A2(n_718), .B(n_719), .Y(n_717) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g822 ( .A(n_641), .Y(n_822) );
INVx2_ASAP7_75t_L g1368 ( .A(n_641), .Y(n_1368) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g690 ( .A(n_642), .Y(n_690) );
INVx1_ASAP7_75t_L g771 ( .A(n_642), .Y(n_771) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx12f_ASAP7_75t_L g676 ( .A(n_647), .Y(n_676) );
BUFx6f_ASAP7_75t_L g1342 ( .A(n_647), .Y(n_1342) );
BUFx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g880 ( .A(n_653), .Y(n_880) );
INVx1_ASAP7_75t_L g1339 ( .A(n_653), .Y(n_1339) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g1349 ( .A(n_663), .Y(n_1349) );
INVx2_ASAP7_75t_L g735 ( .A(n_664), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_705), .B1(n_706), .B2(n_788), .Y(n_666) );
INVx3_ASAP7_75t_L g789 ( .A(n_667), .Y(n_789) );
NAND3xp33_ASAP7_75t_SL g668 ( .A(n_669), .B(n_674), .C(n_681), .Y(n_668) );
BUFx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND3x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .C(n_680), .Y(n_674) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_679), .Y(n_1059) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_691), .C(n_698), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_687), .B2(n_688), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g930 ( .A(n_686), .Y(n_930) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_696), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_757), .B1(n_758), .B2(n_787), .Y(n_707) );
INVx1_ASAP7_75t_L g787 ( .A(n_708), .Y(n_787) );
XNOR2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_736), .Y(n_708) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_711), .B(n_720), .C(n_724), .D(n_730), .Y(n_710) );
NOR2xp67_ASAP7_75t_L g711 ( .A(n_712), .B(n_717), .Y(n_711) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_723), .Y(n_1065) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
BUFx3_ASAP7_75t_L g1337 ( .A(n_728), .Y(n_1337) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_729), .Y(n_1068) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g890 ( .A(n_732), .Y(n_890) );
INVx1_ASAP7_75t_L g923 ( .A(n_732), .Y(n_923) );
INVx2_ASAP7_75t_L g1013 ( .A(n_732), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
XOR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_756), .Y(n_736) );
NOR4xp75_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .C(n_745), .D(n_748), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_746), .B(n_747), .Y(n_745) );
OAI21x1_ASAP7_75t_SL g748 ( .A1(n_749), .A2(n_750), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_753), .Y(n_844) );
INVx2_ASAP7_75t_L g1048 ( .A(n_753), .Y(n_1048) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NAND4xp75_ASAP7_75t_SL g759 ( .A(n_760), .B(n_764), .C(n_769), .D(n_775), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g1335 ( .A(n_762), .Y(n_1335) );
BUFx3_ASAP7_75t_L g1375 ( .A(n_762), .Y(n_1375) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g928 ( .A(n_774), .Y(n_928) );
INVx2_ASAP7_75t_L g1075 ( .A(n_774), .Y(n_1075) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_784), .B2(n_785), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
XNOR2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_916), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_792), .A2(n_793), .B1(n_870), .B2(n_915), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
XNOR2x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_823), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
XNOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_807), .Y(n_798) );
NAND4xp25_ASAP7_75t_L g799 ( .A(n_800), .B(n_804), .C(n_805), .D(n_806), .Y(n_799) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g977 ( .A(n_802), .Y(n_977) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_817), .C(n_820), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .Y(n_809) );
INVx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx4_ASAP7_75t_L g970 ( .A(n_816), .Y(n_970) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_816), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI22x1_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_849), .B1(n_850), .B2(n_869), .Y(n_823) );
INVx2_ASAP7_75t_L g869 ( .A(n_824), .Y(n_869) );
NAND4xp75_ASAP7_75t_L g825 ( .A(n_826), .B(n_830), .C(n_833), .D(n_843), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_838), .Y(n_833) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B(n_837), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g894 ( .A(n_848), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_848), .B(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_848), .B(n_955), .Y(n_954) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_862), .Y(n_851) );
NAND4xp25_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .C(n_856), .D(n_860), .Y(n_852) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_857), .Y(n_1071) );
NAND4xp25_ASAP7_75t_SL g862 ( .A(n_863), .B(n_866), .C(n_867), .D(n_868), .Y(n_862) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
BUFx3_ASAP7_75t_L g915 ( .A(n_871), .Y(n_915) );
OAI22x1_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_910), .B1(n_913), .B2(n_914), .Y(n_871) );
INVx2_ASAP7_75t_L g913 ( .A(n_872), .Y(n_913) );
OA22x2_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_874), .B1(n_895), .B2(n_909), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND4xp75_ASAP7_75t_L g875 ( .A(n_876), .B(n_881), .C(n_886), .D(n_889), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_884), .Y(n_881) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_883), .Y(n_1066) );
AND2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
INVx2_ASAP7_75t_L g909 ( .A(n_895), .Y(n_909) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_902), .Y(n_896) );
NAND4xp25_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .C(n_900), .D(n_901), .Y(n_897) );
NAND4xp25_ASAP7_75t_SL g902 ( .A(n_903), .B(n_906), .C(n_907), .D(n_908), .Y(n_902) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g914 ( .A(n_912), .Y(n_914) );
XNOR2x1_ASAP7_75t_L g916 ( .A(n_917), .B(n_1001), .Y(n_916) );
XNOR2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_959), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_937), .B1(n_957), .B2(n_958), .Y(n_918) );
INVx2_ASAP7_75t_L g958 ( .A(n_919), .Y(n_958) );
OR2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_931), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_927), .C(n_929), .Y(n_921) );
NAND4xp25_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .C(n_934), .D(n_935), .Y(n_931) );
INVx1_ASAP7_75t_L g957 ( .A(n_937), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_939), .A2(n_1134), .B1(n_1136), .B2(n_1137), .Y(n_1133) );
INVx1_ASAP7_75t_L g956 ( .A(n_940), .Y(n_956) );
NAND4xp75_ASAP7_75t_L g940 ( .A(n_941), .B(n_944), .C(n_948), .D(n_951), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
AND2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .Y(n_951) );
AO22x2_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_986), .B2(n_1000), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_972), .C(n_979), .Y(n_963) );
INVx1_ASAP7_75t_L g985 ( .A(n_964), .Y(n_985) );
AND3x2_ASAP7_75t_L g964 ( .A(n_965), .B(n_968), .C(n_971), .Y(n_964) );
INVxp67_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AND4x1_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .C(n_975), .D(n_978), .Y(n_972) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_987), .Y(n_1000) );
NAND3x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .C(n_995), .Y(n_988) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
AND4x1_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .C(n_998), .D(n_999), .Y(n_995) );
AOI21x1_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1054), .B(n_1082), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1003), .B(n_1055), .Y(n_1082) );
OA22x2_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1019), .B1(n_1052), .B2(n_1053), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1004), .Y(n_1052) );
XOR2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1018), .Y(n_1004) );
NOR2x1_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1011), .Y(n_1005) );
NAND4xp25_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .C(n_1009), .D(n_1010), .Y(n_1006) );
NAND4xp25_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1014), .C(n_1015), .D(n_1016), .Y(n_1011) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1019), .Y(n_1053) );
XNOR2x1_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1035), .Y(n_1019) );
XNOR2x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1030), .Y(n_1022) );
NAND4xp25_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .C(n_1026), .D(n_1027), .Y(n_1023) );
NAND4xp25_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1032), .C(n_1033), .D(n_1034), .Y(n_1030) );
XNOR2x1_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1051), .Y(n_1035) );
NAND4xp75_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1040), .C(n_1043), .D(n_1046), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_1055), .Y(n_1054) );
NAND4xp75_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1063), .C(n_1069), .D(n_1076), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1060), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1067), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1073), .Y(n_1069) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1327), .B1(n_1329), .B2(n_1354), .C(n_1358), .Y(n_1083) );
AOI21x1_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1242), .B(n_1291), .Y(n_1084) );
NAND5xp2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1175), .C(n_1205), .D(n_1217), .E(n_1229), .Y(n_1085) );
AOI221xp5_ASAP7_75t_SL g1086 ( .A1(n_1087), .A2(n_1155), .B1(n_1165), .B2(n_1169), .C(n_1170), .Y(n_1086) );
A2O1A1Ixp33_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1139), .B(n_1143), .C(n_1148), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_1088), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1127), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
AOI211xp5_ASAP7_75t_L g1213 ( .A1(n_1090), .A2(n_1206), .B(n_1214), .C(n_1216), .Y(n_1213) );
OAI21xp33_ASAP7_75t_L g1232 ( .A1(n_1090), .A2(n_1233), .B(n_1235), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1113), .Y(n_1090) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1091), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1091), .B(n_1167), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1091), .B(n_1182), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1091), .B(n_1220), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1091), .B(n_1190), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1091), .B(n_1154), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1091), .B(n_1192), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1091), .B(n_1143), .Y(n_1304) );
CKINVDCx6p67_ASAP7_75t_R g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1092), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1092), .B(n_1113), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1092), .B(n_1127), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1092), .B(n_1192), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1092), .B(n_1245), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1092), .B(n_1167), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1092), .B(n_1127), .Y(n_1270) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1092), .B(n_1128), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1092), .B(n_1283), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_1092), .B(n_1268), .Y(n_1288) );
OR2x6_ASAP7_75t_SL g1092 ( .A(n_1093), .B(n_1103), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1099), .B1(n_1100), .B2(n_1102), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1096), .B(n_1101), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_1096), .B(n_1101), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_1096), .B(n_1111), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1096), .B(n_1101), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_1096), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_1100), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_1100), .A2(n_1130), .B1(n_1201), .B2(n_1202), .C(n_1203), .Y(n_1200) );
BUFx2_ASAP7_75t_L g1328 ( .A(n_1100), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1101), .B(n_1107), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1101), .B(n_1107), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1101), .B(n_1107), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_1104), .A2(n_1105), .B1(n_1108), .B2(n_1109), .Y(n_1103) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1107), .B(n_1111), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1107), .B(n_1111), .Y(n_1122) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1107), .B(n_1111), .Y(n_1135) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1113), .B(n_1140), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1113), .B(n_1167), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1113), .B(n_1210), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1113), .B(n_1193), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1119), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1114), .B(n_1140), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1114), .B(n_1120), .Y(n_1174) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_1115), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1115), .B(n_1120), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1115), .B(n_1119), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1115), .B(n_1140), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1115), .B(n_1140), .Y(n_1299) );
AND2x4_ASAP7_75t_SL g1115 ( .A(n_1116), .B(n_1118), .Y(n_1115) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1117), .Y(n_1164) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1119), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1119), .B(n_1182), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1119), .B(n_1182), .Y(n_1283) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1124), .Y(n_1120) );
INVx3_ASAP7_75t_L g1130 ( .A(n_1125), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1127), .B(n_1145), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1127), .B(n_1184), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1127), .B(n_1159), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1127), .B(n_1158), .Y(n_1250) );
INVx3_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1128), .B(n_1144), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1128), .B(n_1145), .Y(n_1190) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1128), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1128), .B(n_1145), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1133), .Y(n_1128) );
INVx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1139), .Y(n_1321) );
CKINVDCx6p67_ASAP7_75t_R g1167 ( .A(n_1140), .Y(n_1167) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1140), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1140), .B(n_1221), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1140), .B(n_1174), .Y(n_1245) );
OAI322xp33_ASAP7_75t_L g1251 ( .A1(n_1140), .A2(n_1157), .A3(n_1252), .B1(n_1253), .B2(n_1256), .C1(n_1257), .C2(n_1259), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_1143), .A2(n_1230), .B1(n_1231), .B2(n_1232), .C(n_1236), .Y(n_1229) );
INVx3_ASAP7_75t_L g1271 ( .A(n_1143), .Y(n_1271) );
OAI21xp5_ASAP7_75t_L g1272 ( .A1(n_1143), .A2(n_1273), .B(n_1274), .Y(n_1272) );
INVx3_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1144), .B(n_1160), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1144), .B(n_1160), .Y(n_1195) );
INVx2_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1145), .B(n_1160), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1149), .B(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1151), .B(n_1180), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1151), .B(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1154), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1152), .B(n_1174), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1152), .B(n_1160), .Y(n_1287) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1152), .B(n_1317), .Y(n_1316) );
O2A1O1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1152), .A2(n_1187), .B(n_1196), .C(n_1240), .Y(n_1326) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1154), .B(n_1157), .Y(n_1280) );
NAND3xp33_ASAP7_75t_L g1323 ( .A(n_1154), .B(n_1226), .C(n_1287), .Y(n_1323) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1155), .Y(n_1309) );
INVx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx3_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1157), .B(n_1171), .Y(n_1170) );
INVx3_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1159), .B(n_1198), .Y(n_1197) );
A2O1A1Ixp33_ASAP7_75t_L g1320 ( .A1(n_1159), .A2(n_1189), .B(n_1321), .C(n_1322), .Y(n_1320) );
INVx3_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1160), .B(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1160), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1160), .B(n_1264), .Y(n_1296) );
AND2x4_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .Y(n_1166) );
AND2x2_ASAP7_75t_SL g1173 ( .A(n_1167), .B(n_1174), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_1167), .B(n_1212), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1167), .B(n_1221), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1167), .B(n_1192), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1168), .B(n_1182), .Y(n_1273) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1168), .Y(n_1298) );
AOI322xp5_ASAP7_75t_L g1294 ( .A1(n_1169), .A2(n_1218), .A3(n_1258), .B1(n_1295), .B2(n_1297), .C1(n_1299), .C2(n_1300), .Y(n_1294) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_1171), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1239 ( .A(n_1172), .Y(n_1239) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1173), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1174), .B(n_1193), .Y(n_1198) );
AOI222xp33_ASAP7_75t_L g1217 ( .A1(n_1174), .A2(n_1218), .B1(n_1222), .B2(n_1223), .C1(n_1224), .C2(n_1228), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1174), .B(n_1221), .Y(n_1286) );
INVxp33_ASAP7_75t_L g1317 ( .A(n_1174), .Y(n_1317) );
NOR3xp33_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1194), .C(n_1204), .Y(n_1175) );
OAI32xp33_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1184), .A3(n_1185), .B1(n_1187), .B2(n_1191), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1179), .Y(n_1278) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1180), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
AOI321xp33_ASAP7_75t_L g1285 ( .A1(n_1182), .A2(n_1231), .A3(n_1286), .B1(n_1287), .B2(n_1288), .C(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1184), .Y(n_1222) );
OAI211xp5_ASAP7_75t_L g1319 ( .A1(n_1184), .A2(n_1275), .B(n_1320), .C(n_1323), .Y(n_1319) );
CKINVDCx14_ASAP7_75t_R g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1262 ( .A1(n_1190), .A2(n_1263), .B1(n_1265), .B2(n_1266), .C(n_1269), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1192), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1192), .B(n_1247), .Y(n_1246) );
NAND3xp33_ASAP7_75t_L g1269 ( .A(n_1192), .B(n_1270), .C(n_1271), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1192), .B(n_1210), .Y(n_1308) );
OAI211xp5_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1196), .B(n_1197), .C(n_1199), .Y(n_1194) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1195), .Y(n_1216) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1197), .Y(n_1322) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1200), .Y(n_1290) );
AOI211xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1209), .B(n_1211), .C(n_1213), .Y(n_1205) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1208), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1208), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1209), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1214), .B(n_1253), .Y(n_1284) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1216), .B(n_1234), .Y(n_1258) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_1216), .A2(n_1278), .B1(n_1279), .B2(n_1281), .C(n_1284), .Y(n_1277) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1221), .Y(n_1268) );
AOI21xp5_ASAP7_75t_L g1260 ( .A1(n_1222), .A2(n_1261), .B(n_1262), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1227), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1228), .Y(n_1318) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1234), .B(n_1308), .Y(n_1307) );
AOI21xp5_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1239), .B(n_1240), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
O2A1O1Ixp33_ASAP7_75t_L g1324 ( .A1(n_1238), .A2(n_1246), .B(n_1325), .C(n_1326), .Y(n_1324) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NAND5xp2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1260), .C(n_1272), .D(n_1277), .E(n_1285), .Y(n_1242) );
O2A1O1Ixp33_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1246), .B(n_1249), .C(n_1251), .Y(n_1243) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1245), .Y(n_1314) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1246), .Y(n_1265) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1248), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_SL g1297 ( .A(n_1248), .B(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVxp67_ASAP7_75t_SL g1274 ( .A(n_1275), .Y(n_1274) );
AOI21xp33_ASAP7_75t_L g1310 ( .A1(n_1279), .A2(n_1311), .B(n_1313), .Y(n_1310) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1324), .Y(n_1291) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1319), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1302), .C(n_1310), .Y(n_1293) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
A2O1A1Ixp33_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1305), .B(n_1306), .C(n_1309), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
AOI21xp33_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1315), .B(n_1318), .Y(n_1313) );
INVxp33_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1343), .Y(n_1331) );
NAND4xp25_ASAP7_75t_SL g1332 ( .A(n_1333), .B(n_1336), .C(n_1338), .D(n_1341), .Y(n_1332) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1351), .C(n_1353), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
OAI21xp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B(n_1350), .Y(n_1347) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVxp67_ASAP7_75t_SL g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
NOR2x1_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1371), .Y(n_1363) );
NAND4xp25_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1367), .C(n_1369), .D(n_1370), .Y(n_1364) );
NAND4xp25_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1374), .C(n_1376), .D(n_1377), .Y(n_1371) );
BUFx3_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
endmodule