module fake_jpeg_18931_n_288 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_29),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_57),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_33),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_26),
.B(n_16),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_101),
.B(n_30),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_96),
.B1(n_97),
.B2(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_66),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_18),
.B1(n_14),
.B2(n_24),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_16),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_18),
.B1(n_24),
.B2(n_37),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_35),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_39),
.B1(n_41),
.B2(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_39),
.B1(n_44),
.B2(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_44),
.B1(n_42),
.B2(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_15),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_32),
.B1(n_31),
.B2(n_34),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_87),
.B1(n_32),
.B2(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_19),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_26),
.B1(n_30),
.B2(n_23),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_100),
.B1(n_91),
.B2(n_81),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_35),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_43),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_21),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_43),
.B(n_1),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_29),
.B(n_17),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_124),
.B(n_132),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_121),
.B1(n_96),
.B2(n_20),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_31),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_22),
.A3(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_67),
.B(n_96),
.C(n_17),
.D(n_77),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_69),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_70),
.B(n_17),
.Y(n_132)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_75),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_148),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_115),
.B1(n_122),
.B2(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_61),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_61),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_147),
.Y(n_175)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_100),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_79),
.B(n_78),
.C(n_82),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_155),
.B(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_62),
.B1(n_76),
.B2(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_114),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_108),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_93),
.B1(n_17),
.B2(n_98),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_111),
.B1(n_128),
.B2(n_129),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_84),
.B1(n_8),
.B2(n_13),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_88),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_145),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_113),
.C(n_109),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_153),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_168),
.B1(n_160),
.B2(n_154),
.Y(n_200)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_124),
.B(n_130),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_144),
.B(n_142),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_185),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_116),
.B1(n_128),
.B2(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_186),
.B1(n_158),
.B2(n_148),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_106),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_129),
.B1(n_117),
.B2(n_126),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_7),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_149),
.B(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_144),
.B(n_155),
.C(n_147),
.D(n_134),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_194),
.B(n_195),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_147),
.B(n_150),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_210),
.B1(n_170),
.B2(n_177),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_120),
.B(n_108),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_184),
.B(n_161),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_206),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_171),
.B(n_182),
.C(n_164),
.D(n_174),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_135),
.B(n_85),
.C(n_104),
.D(n_8),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_184),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_162),
.B(n_11),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_104),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_186),
.C(n_173),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_161),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_141),
.B1(n_10),
.B2(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_199),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_216),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_230),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_187),
.C(n_163),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_229),
.C(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_227),
.B1(n_228),
.B2(n_181),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_201),
.B(n_197),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_141),
.C(n_169),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_172),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_198),
.C(n_203),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_188),
.B1(n_192),
.B2(n_207),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_236),
.B1(n_232),
.B2(n_240),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_188),
.B(n_207),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_240),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_188),
.CI(n_210),
.CON(n_239),
.SN(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_188),
.C(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_172),
.C(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_181),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_215),
.C(n_230),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_167),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_227),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_218),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_216),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_235),
.B(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_264),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_259),
.A2(n_242),
.B(n_233),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_267),
.B(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_243),
.C(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_245),
.B(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_270),
.A3(n_263),
.B1(n_260),
.B2(n_179),
.C1(n_3),
.C2(n_4),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_248),
.C(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.C(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_247),
.C(n_239),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_239),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_279),
.C(n_179),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_179),
.B(n_1),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_0),
.B(n_2),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_283),
.A3(n_282),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_0),
.C(n_2),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_3),
.C(n_4),
.Y(n_288)
);


endmodule