module fake_jpeg_32111_n_185 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_52),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_71),
.B1(n_69),
.B2(n_76),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_64),
.B(n_67),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_61),
.B1(n_69),
.B2(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_71),
.B1(n_76),
.B2(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_72),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_78),
.CI(n_82),
.CON(n_108),
.SN(n_108)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_51),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_84),
.B1(n_81),
.B2(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_91),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_67),
.C(n_66),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_0),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_7),
.Y(n_141)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_75),
.B1(n_70),
.B2(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_77),
.B1(n_74),
.B2(n_68),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_129),
.B(n_140),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_22),
.B1(n_50),
.B2(n_48),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_19),
.B(n_45),
.C(n_43),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_138),
.B1(n_9),
.B2(n_10),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_18),
.B1(n_41),
.B2(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_4),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_122),
.C(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_157),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_119),
.A3(n_101),
.B1(n_24),
.B2(n_27),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_106),
.C(n_39),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_38),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_120),
.B(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_8),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_8),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_152),
.C(n_149),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_164),
.B1(n_156),
.B2(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_172),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_161),
.A3(n_176),
.B1(n_168),
.B2(n_170),
.C1(n_154),
.C2(n_163),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_167),
.B(n_143),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_147),
.B(n_165),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_23),
.A3(n_34),
.B1(n_32),
.B2(n_29),
.C1(n_155),
.C2(n_16),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_15),
.C(n_16),
.Y(n_185)
);


endmodule