module real_aes_6711_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_10;
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_0), .B(n_4), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_2), .B(n_14), .Y(n_13) );
CKINVDCx14_ASAP7_75t_R g25 ( .A(n_2), .Y(n_25) );
NAND3xp33_ASAP7_75t_SL g10 ( .A(n_3), .B(n_11), .C(n_12), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_4), .B(n_21), .Y(n_20) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g27 ( .A(n_6), .Y(n_27) );
INVx2_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
AOI21xp33_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_15), .B(n_23), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx1_ASAP7_75t_SL g12 ( .A(n_13), .Y(n_12) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_14), .B(n_25), .C(n_26), .Y(n_24) );
OAI22xp33_ASAP7_75t_L g15 ( .A1(n_16), .A2(n_17), .B1(n_20), .B2(n_22), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_24), .Y(n_23) );
INVx1_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
endmodule