module fake_jpeg_24825_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_15),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_23),
.B(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_71),
.Y(n_89)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_86),
.B1(n_54),
.B2(n_23),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_70),
.B1(n_77),
.B2(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_26),
.B1(n_31),
.B2(n_21),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_66),
.B1(n_19),
.B2(n_30),
.Y(n_107)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_0),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_69),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_24),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_73),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_83),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_30),
.B1(n_24),
.B2(n_27),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_53),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_29),
.B1(n_16),
.B2(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_79),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_111),
.B(n_63),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_107),
.B1(n_65),
.B2(n_85),
.Y(n_120)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_65),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_55),
.A3(n_25),
.B1(n_30),
.B2(n_53),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_80),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_30),
.B1(n_53),
.B2(n_24),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_24),
.C(n_1),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_70),
.C(n_83),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_76),
.B1(n_60),
.B2(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_124),
.B1(n_57),
.B2(n_62),
.Y(n_168)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_57),
.B1(n_62),
.B2(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_129),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_95),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_140),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_15),
.B(n_14),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_74),
.C(n_64),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_101),
.C(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_64),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_79),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_115),
.B(n_138),
.C(n_139),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_143),
.B(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_160),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_111),
.B(n_110),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_87),
.B(n_111),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_87),
.B1(n_91),
.B2(n_105),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_152),
.B1(n_162),
.B2(n_129),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_109),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_165),
.C(n_166),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_164),
.B(n_84),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_157),
.Y(n_172)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_8),
.B(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_81),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_170),
.B(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_136),
.B1(n_140),
.B2(n_116),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_67),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_97),
.C(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_116),
.B(n_123),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_96),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_14),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_98),
.B(n_84),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_180),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_124),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_122),
.C(n_118),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_118),
.B1(n_117),
.B2(n_128),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_127),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_117),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_164),
.B(n_145),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_191),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_1),
.B(n_2),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_143),
.B(n_146),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_119),
.C(n_112),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_188),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_207),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_164),
.B(n_169),
.C(n_147),
.D(n_151),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_193),
.C(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_197),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_149),
.B1(n_167),
.B2(n_146),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_214),
.B1(n_175),
.B2(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_154),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_181),
.B1(n_171),
.B2(n_149),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_173),
.B(n_174),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_225),
.B(n_226),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_229),
.B(n_203),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_227),
.B1(n_207),
.B2(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_171),
.B1(n_192),
.B2(n_155),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_183),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_205),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_199),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_237),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_200),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_229),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_215),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_228),
.C(n_204),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_158),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_252),
.C(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_217),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

AOI31xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_221),
.A3(n_242),
.B(n_241),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_253),
.B(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_230),
.B1(n_209),
.B2(n_224),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_161),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_161),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_208),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_249),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_157),
.B1(n_195),
.B2(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_261),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_10),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_14),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_266),
.C(n_271),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_253),
.A3(n_249),
.B1(n_252),
.B2(n_12),
.C1(n_7),
.C2(n_11),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_258),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_7),
.B(n_12),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_11),
.B(n_13),
.C(n_5),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_265),
.B(n_267),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_278),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_4),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_4),
.B(n_5),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_274),
.C1(n_250),
.C2(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_274),
.C(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_6),
.Y(n_283)
);


endmodule