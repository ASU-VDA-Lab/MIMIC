module fake_jpeg_16246_n_156 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_156);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_5),
.B(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_5),
.B(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_34),
.B(n_36),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_41),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_48),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_5),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_28),
.B1(n_18),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_70),
.B1(n_60),
.B2(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_13),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_28),
.B1(n_15),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_60),
.B1(n_51),
.B2(n_59),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_8),
.B(n_12),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_14),
.B1(n_15),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_14),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_40),
.B(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_19),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_90),
.B1(n_66),
.B2(n_52),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_81),
.B(n_88),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_R g81 ( 
.A(n_55),
.B(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_40),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_97),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_8),
.B1(n_12),
.B2(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_71),
.B1(n_52),
.B2(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_71),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_106),
.B1(n_110),
.B2(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_85),
.B1(n_94),
.B2(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_72),
.B1(n_53),
.B2(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_53),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_89),
.C(n_88),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_122),
.C(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_93),
.B1(n_95),
.B2(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_80),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_116),
.B(n_99),
.Y(n_131)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_113),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_105),
.B(n_112),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_80),
.B1(n_92),
.B2(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_134),
.C(n_137),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_118),
.B1(n_129),
.B2(n_127),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_113),
.C(n_103),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_101),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_132),
.C(n_134),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_121),
.A3(n_128),
.B1(n_126),
.B2(n_124),
.C(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

AO221x1_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_125),
.B1(n_111),
.B2(n_112),
.C(n_105),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_149),
.B(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_126),
.Y(n_151)
);

OAI31xp33_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_152),
.A3(n_144),
.B(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_139),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_154),
.Y(n_156)
);


endmodule