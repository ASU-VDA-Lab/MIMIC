module real_jpeg_25360_n_20 (n_17, n_8, n_0, n_93, n_2, n_10, n_9, n_12, n_92, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_94, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_93;
input n_2;
input n_10;
input n_9;
input n_12;
input n_92;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_94;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_50),
.B1(n_57),
.B2(n_68),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_0),
.B(n_76),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_8),
.B1(n_32),
.B2(n_39),
.C(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_3),
.B(n_92),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_94),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_6),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_9),
.B1(n_32),
.B2(n_41),
.C(n_42),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_15),
.B1(n_32),
.B2(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_11),
.B1(n_32),
.B2(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_47),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_17),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_13),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_93),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_22),
.B1(n_23),
.B2(n_48),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_19),
.A2(n_48),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_49),
.B1(n_75),
.B2(n_79),
.C(n_89),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR5xp2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.C(n_44),
.D(n_45),
.E(n_47),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_26),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_32),
.C(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR5xp2_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_38),
.C(n_45),
.D(n_82),
.E(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_59),
.B(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_70),
.B(n_73),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_73),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_64),
.B(n_67),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_88),
.Y(n_87)
);


endmodule