module fake_jpeg_26648_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_28),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_18),
.B1(n_16),
.B2(n_30),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_55),
.B1(n_17),
.B2(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_16),
.B1(n_30),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_62),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_26),
.B1(n_27),
.B2(n_22),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_58),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_51),
.B(n_54),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_21),
.C(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_88),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_22),
.B(n_25),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_27),
.B(n_25),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_31),
.B1(n_24),
.B2(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_91),
.B1(n_64),
.B2(n_60),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_20),
.B1(n_24),
.B2(n_17),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_33),
.B(n_29),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_33),
.B1(n_20),
.B2(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_44),
.A2(n_19),
.B1(n_29),
.B2(n_20),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_45),
.B1(n_57),
.B2(n_33),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_101),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_61),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_46),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_116),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_66),
.B1(n_69),
.B2(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_77),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_85),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_135),
.B(n_140),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_69),
.C(n_68),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_126),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_87),
.B1(n_77),
.B2(n_84),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_125),
.B1(n_131),
.B2(n_139),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_128),
.Y(n_154)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_133),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_84),
.B1(n_83),
.B2(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_136),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_138),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_83),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_74),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_90),
.B1(n_72),
.B2(n_73),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_155),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_107),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_92),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_109),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_94),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_116),
.B1(n_113),
.B2(n_106),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_123),
.B1(n_139),
.B2(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_89),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_99),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_192),
.B1(n_189),
.B2(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_160),
.B1(n_151),
.B2(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_118),
.B1(n_140),
.B2(n_127),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_143),
.C(n_109),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_168),
.C(n_170),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_144),
.B1(n_111),
.B2(n_78),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_144),
.B1(n_111),
.B2(n_78),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_197),
.B1(n_152),
.B2(n_143),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_80),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_76),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_81),
.B1(n_100),
.B2(n_33),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_148),
.B1(n_146),
.B2(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_221),
.B1(n_193),
.B2(n_176),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_215),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_205),
.B1(n_208),
.B2(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_186),
.B1(n_196),
.B2(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_149),
.B1(n_164),
.B2(n_163),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_218),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_213),
.C(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_158),
.C(n_145),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_171),
.B(n_158),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_169),
.C(n_145),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_70),
.B1(n_60),
.B2(n_52),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_70),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_208),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_234),
.B1(n_224),
.B2(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_184),
.B1(n_181),
.B2(n_188),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_185),
.C(n_70),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_52),
.C(n_8),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_213),
.B1(n_206),
.B2(n_214),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_219),
.B(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_217),
.B1(n_204),
.B2(n_3),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_248),
.B1(n_253),
.B2(n_229),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_217),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_233),
.C(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_223),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_7),
.B(n_14),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_235),
.B(n_15),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_265),
.B1(n_10),
.B2(n_15),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_228),
.B1(n_238),
.B2(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_223),
.C(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_251),
.Y(n_271)
);

AOI211xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_10),
.B(n_14),
.C(n_5),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_244),
.B(n_242),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_257),
.B1(n_264),
.B2(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_272),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_252),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_265),
.A3(n_260),
.B1(n_6),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_275),
.C(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_263),
.B(n_6),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_12),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_6),
.B(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_275),
.B(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_276),
.C(n_281),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_287),
.B(n_285),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_289),
.C(n_286),
.Y(n_291)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_1),
.A3(n_4),
.B1(n_15),
.B2(n_277),
.C(n_290),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_1),
.Y(n_293)
);


endmodule