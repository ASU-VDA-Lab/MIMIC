module fake_jpeg_5323_n_109 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_24),
.B1(n_8),
.B2(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_8),
.B1(n_21),
.B2(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_28),
.B1(n_13),
.B2(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_19),
.B(n_20),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_12),
.B(n_11),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_46),
.B1(n_18),
.B2(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_26),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_33),
.B1(n_41),
.B2(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_38),
.C(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_42),
.C(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_12),
.C(n_3),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_43),
.B(n_50),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_75),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_43),
.B(n_12),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_62),
.B(n_65),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.C(n_64),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_37),
.C(n_18),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_17),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AO221x1_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_75),
.B1(n_68),
.B2(n_80),
.C(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_58),
.C(n_54),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_76),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_96),
.B1(n_37),
.B2(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_58),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_84),
.B1(n_17),
.B2(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_91),
.B1(n_77),
.B2(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_6),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_0),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_48),
.C2(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_100),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_103),
.B(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_7),
.Y(n_109)
);


endmodule