module fake_jpeg_29819_n_418 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_17),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_60),
.Y(n_89)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_71),
.Y(n_102)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_0),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_32),
.B(n_16),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_79),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_26),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_41),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_34),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_85),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_97),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_133),
.B1(n_136),
.B2(n_22),
.Y(n_148)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_34),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_48),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_70),
.B(n_41),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_105),
.Y(n_140)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_46),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_52),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_38),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_158),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_58),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_151),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_163),
.B1(n_88),
.B2(n_117),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_94),
.A2(n_36),
.B1(n_47),
.B2(n_53),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_107),
.B1(n_124),
.B2(n_96),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_101),
.C(n_116),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_38),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_157),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_109),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_95),
.B(n_49),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_171),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_86),
.B(n_18),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_165),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_92),
.A2(n_59),
.B1(n_69),
.B2(n_54),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_79),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_108),
.A2(n_36),
.B1(n_75),
.B2(n_68),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_92),
.A2(n_57),
.B1(n_62),
.B2(n_61),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_135),
.B1(n_100),
.B2(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_104),
.B1(n_100),
.B2(n_106),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_179),
.B1(n_173),
.B2(n_175),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_132),
.B(n_123),
.C(n_111),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_187),
.B(n_145),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_88),
.B1(n_106),
.B2(n_117),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_142),
.B1(n_171),
.B2(n_167),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_111),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_132),
.B(n_110),
.C(n_103),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_144),
.B(n_166),
.C(n_153),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_194),
.B1(n_200),
.B2(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_181),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_204),
.Y(n_219)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_173),
.B1(n_185),
.B2(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_143),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_174),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_167),
.B(n_107),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_209),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_212),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_158),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_191),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_197),
.B(n_206),
.Y(n_234)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_152),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_200),
.B1(n_204),
.B2(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_220),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_197),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_178),
.B1(n_173),
.B2(n_179),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_225),
.B1(n_194),
.B2(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_231),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_174),
.A3(n_187),
.B1(n_186),
.B2(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_142),
.B1(n_193),
.B2(n_155),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_205),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_192),
.B(n_190),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_190),
.A3(n_182),
.B1(n_161),
.B2(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_206),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_218),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_196),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_253),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_213),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_214),
.B(n_209),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_207),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_223),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_218),
.C(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_251),
.C(n_244),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_223),
.Y(n_260)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_262),
.Y(n_283)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_214),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_264),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_228),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_265),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_237),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_226),
.B(n_229),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_229),
.B(n_236),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_219),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_249),
.B1(n_220),
.B2(n_216),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_245),
.C(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_259),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_255),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_235),
.B1(n_236),
.B2(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_291),
.B1(n_265),
.B2(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_295),
.B1(n_298),
.B2(n_225),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_224),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_293),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_264),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_230),
.B1(n_224),
.B2(n_237),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_203),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_274),
.Y(n_321)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_229),
.B1(n_205),
.B2(n_240),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_300),
.B1(n_202),
.B2(n_208),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_294),
.A2(n_256),
.B1(n_289),
.B2(n_282),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_298),
.C(n_231),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_271),
.CI(n_255),
.CON(n_304),
.SN(n_304)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_315),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_276),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_307),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_287),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_272),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_306),
.C(n_305),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_284),
.A2(n_263),
.B1(n_269),
.B2(n_266),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_318),
.B1(n_322),
.B2(n_208),
.Y(n_334)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_273),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_211),
.Y(n_340)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_284),
.A2(n_266),
.B1(n_257),
.B2(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_320),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_321),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_257),
.B1(n_261),
.B2(n_239),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_334),
.Y(n_360)
);

A2O1A1O1Ixp25_ASAP7_75t_L g325 ( 
.A1(n_301),
.A2(n_261),
.B(n_227),
.C(n_209),
.D(n_283),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_152),
.C(n_169),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_311),
.A2(n_290),
.B(n_283),
.C(n_295),
.Y(n_327)
);

AOI21x1_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_338),
.B(n_137),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_160),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_232),
.C(n_203),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_330),
.B(n_332),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_331),
.A2(n_339),
.B1(n_141),
.B2(n_113),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_180),
.C(n_182),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_202),
.B(n_208),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_302),
.A2(n_202),
.B1(n_211),
.B2(n_142),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_316),
.Y(n_346)
);

INVx13_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_211),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_152),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_310),
.B1(n_312),
.B2(n_309),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_345),
.A2(n_325),
.B1(n_327),
.B2(n_342),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_349),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_322),
.B(n_180),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_347),
.A2(n_356),
.B(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_350),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_344),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_354),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_180),
.C(n_169),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_355),
.C(n_358),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_353),
.B(n_340),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_160),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_137),
.C(n_154),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_164),
.B(n_141),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_357),
.A2(n_335),
.B1(n_343),
.B2(n_328),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_137),
.C(n_115),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_93),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_336),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_366),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_112),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_370),
.B1(n_376),
.B2(n_350),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_362),
.A2(n_327),
.B1(n_338),
.B2(n_36),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_371),
.B(n_372),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_96),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_372),
.A2(n_375),
.B1(n_125),
.B2(n_118),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_112),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_124),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_348),
.A2(n_115),
.B1(n_99),
.B2(n_121),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_381),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_368),
.A2(n_360),
.B1(n_355),
.B2(n_354),
.Y(n_378)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

AOI321xp33_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_360),
.A3(n_358),
.B1(n_346),
.B2(n_110),
.C(n_103),
.Y(n_379)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_375),
.B(n_364),
.Y(n_380)
);

XNOR2x2_ASAP7_75t_SL g389 ( 
.A(n_380),
.B(n_385),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_369),
.B(n_13),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_386),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_14),
.B(n_12),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_369),
.B(n_12),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_388),
.C(n_386),
.Y(n_394)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_373),
.A3(n_28),
.B1(n_131),
.B2(n_77),
.C1(n_42),
.C2(n_14),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_391),
.A2(n_10),
.B(n_22),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_392),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_125),
.C(n_118),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_395),
.A2(n_396),
.B(n_398),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_14),
.C(n_10),
.Y(n_396)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g408 ( 
.A1(n_400),
.A2(n_401),
.A3(n_405),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_22),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_402),
.B(n_403),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_397),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_404),
.A2(n_1),
.B(n_2),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

OAI21xp33_ASAP7_75t_L g406 ( 
.A1(n_399),
.A2(n_389),
.B(n_391),
.Y(n_406)
);

AOI31xp33_ASAP7_75t_L g412 ( 
.A1(n_406),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_SL g413 ( 
.A1(n_408),
.A2(n_407),
.B(n_5),
.C(n_6),
.Y(n_413)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_1),
.B(n_2),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_4),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_413),
.B1(n_409),
.B2(n_29),
.Y(n_414)
);

AOI322xp5_ASAP7_75t_SL g416 ( 
.A1(n_414),
.A2(n_415),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_29),
.C2(n_152),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_6),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_417),
.B(n_7),
.Y(n_418)
);


endmodule