module fake_netlist_6_1150_n_1676 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1676);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1676;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_87),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_14),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_40),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_49),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_68),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_69),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_13),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_54),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_129),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_17),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_64),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_40),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_43),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_103),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_74),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_42),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_104),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_18),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_4),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_31),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_21),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_72),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_31),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_49),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_44),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_63),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_58),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_95),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_98),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_79),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_146),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_73),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_13),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_81),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_57),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_30),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_139),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_102),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_28),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_54),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_77),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_110),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_17),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_5),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_44),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_52),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_26),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_96),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_11),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_90),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_114),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_21),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_59),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_94),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_155),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_29),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_86),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_147),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

INVx4_ASAP7_75t_R g300 ( 
.A(n_158),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_10),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_23),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_109),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_45),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_141),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_34),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_144),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_71),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_47),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_36),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_62),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_170),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_170),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_228),
.B(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_170),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_228),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_229),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_213),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_171),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_213),
.Y(n_323)
);

BUFx2_ASAP7_75t_SL g324 ( 
.A(n_181),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_2),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_167),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_213),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_213),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_213),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_168),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_194),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_197),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_172),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_173),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_187),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_171),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_178),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_185),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_207),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_171),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_190),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_180),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_2),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_192),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_193),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_251),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_312),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_259),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_272),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_272),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_200),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_174),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_202),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_204),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_161),
.B(n_3),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_231),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_161),
.B(n_175),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_175),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_206),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_231),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_174),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_210),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_217),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_222),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_183),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_183),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_312),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_195),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_160),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

BUFx12f_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_191),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_387),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_232),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_229),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_233),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_376),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_235),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_322),
.B(n_244),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

AND3x2_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_220),
.C(n_191),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_324),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_331),
.B(n_236),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_331),
.B(n_238),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_241),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_245),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_244),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_319),
.B(n_306),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

XNOR2x2_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_209),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_246),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_357),
.B(n_306),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_358),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_327),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_252),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_386),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_423),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_333),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_391),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_391),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_397),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_340),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

AND3x2_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_216),
.C(n_179),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_408),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_337),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_431),
.B(n_338),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_415),
.B(n_343),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_344),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_449),
.A2(n_225),
.B1(n_294),
.B2(n_302),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_389),
.B(n_354),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_408),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_422),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_400),
.B(n_347),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_359),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_437),
.B(n_186),
.C(n_184),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_426),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_426),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_400),
.B(n_348),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_374),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_394),
.B(n_184),
.Y(n_507)
);

BUFx6f_ASAP7_75t_SL g508 ( 
.A(n_455),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_409),
.B(n_355),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_409),
.B(n_356),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_398),
.B(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_392),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_398),
.B(n_372),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_388),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_434),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_401),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_417),
.A2(n_254),
.B1(n_240),
.B2(n_224),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_427),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_395),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_434),
.B(n_377),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_438),
.B(n_220),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_437),
.B(n_381),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_417),
.A2(n_212),
.B1(n_288),
.B2(n_378),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_255),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_417),
.A2(n_254),
.B1(n_224),
.B2(n_240),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_428),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_455),
.B(n_371),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_417),
.A2(n_242),
.B1(n_269),
.B2(n_195),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_450),
.B(n_258),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_402),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_457),
.B(n_260),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_401),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_401),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_441),
.A2(n_394),
.B1(n_449),
.B2(n_457),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_441),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_403),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_401),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_455),
.B(n_382),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_449),
.B(n_334),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_389),
.B(n_380),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_394),
.B(n_188),
.C(n_186),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_403),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_424),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_405),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_389),
.B(n_176),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_410),
.B(n_268),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_402),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_412),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_419),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_394),
.A2(n_198),
.B1(n_242),
.B2(n_302),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_453),
.B(n_176),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g573 ( 
.A(n_453),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_419),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_394),
.A2(n_269),
.B1(n_278),
.B2(n_294),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_413),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_414),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_410),
.B(n_270),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_453),
.B(n_182),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_414),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_416),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_416),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_410),
.B(n_271),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_410),
.B(n_182),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_424),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_420),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_439),
.B(n_324),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_439),
.B(n_440),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_421),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_402),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_425),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_425),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_430),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_410),
.A2(n_211),
.B1(n_248),
.B2(n_265),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_440),
.A2(n_278),
.B1(n_296),
.B2(n_208),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_430),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_424),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_444),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_444),
.B(n_182),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_447),
.B(n_176),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_433),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_411),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_411),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_463),
.B(n_283),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_498),
.B(n_499),
.Y(n_608)
);

BUFx5_ASAP7_75t_L g609 ( 
.A(n_584),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_464),
.B(n_447),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_524),
.B(n_402),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_335),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_553),
.A2(n_361),
.B1(n_345),
.B2(n_166),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_SL g614 ( 
.A(n_596),
.B(n_280),
.C(n_277),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_520),
.B(n_490),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_480),
.A2(n_296),
.B1(n_188),
.B2(n_201),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_475),
.B(n_404),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_474),
.A2(n_411),
.B(n_205),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_553),
.B(n_182),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_514),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_476),
.B(n_470),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_470),
.B(n_182),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_492),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_486),
.B(n_163),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_481),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_486),
.B(n_404),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_589),
.A2(n_461),
.B(n_460),
.C(n_458),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_501),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_567),
.A2(n_436),
.B(n_433),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_514),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_487),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_487),
.B(n_201),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_500),
.B(n_404),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_509),
.B(n_404),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_472),
.B(n_164),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_570),
.B(n_205),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_526),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_530),
.B(n_404),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_488),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_589),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_588),
.B(n_279),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_165),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_552),
.B(n_284),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_464),
.B(n_465),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_492),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_462),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_489),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_584),
.B(n_404),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_570),
.A2(n_461),
.B(n_460),
.C(n_458),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_484),
.B(n_176),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_584),
.B(n_436),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

BUFx12f_ASAP7_75t_SL g656 ( 
.A(n_507),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_478),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_572),
.A2(n_237),
.B(n_250),
.C(n_249),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_478),
.Y(n_660)
);

INVx8_ASAP7_75t_L g661 ( 
.A(n_508),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_545),
.B(n_456),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_508),
.A2(n_303),
.B1(n_305),
.B2(n_309),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_531),
.B(n_196),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_496),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_548),
.B(n_456),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_483),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_480),
.A2(n_223),
.B1(n_230),
.B2(n_234),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_483),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_505),
.B(n_169),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_473),
.B(n_177),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_485),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_496),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_502),
.B(n_456),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_502),
.B(n_456),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_531),
.B(n_196),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_513),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_513),
.B(n_519),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_519),
.B(n_411),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_525),
.B(n_411),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_199),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_459),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_529),
.B(n_533),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_529),
.B(n_459),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_534),
.B(n_223),
.C(n_221),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_543),
.B(n_443),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_542),
.B(n_196),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_485),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_479),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_543),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_555),
.B(n_443),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_512),
.B(n_214),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_562),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_515),
.B(n_215),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_542),
.B(n_196),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_562),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_508),
.A2(n_293),
.B1(n_208),
.B2(n_218),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_578),
.A2(n_230),
.B(n_221),
.Y(n_699)
);

BUFx5_ASAP7_75t_L g700 ( 
.A(n_501),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_484),
.B(n_203),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_540),
.B(n_442),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_466),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_462),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_564),
.B(n_459),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_494),
.A2(n_243),
.B(n_295),
.C(n_293),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_484),
.B(n_522),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_574),
.B(n_218),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_484),
.B(n_231),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_542),
.B(n_297),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_542),
.B(n_297),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_507),
.B(n_219),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_494),
.A2(n_507),
.B(n_595),
.C(n_603),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_467),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_467),
.B(n_231),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_577),
.B(n_443),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_580),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_536),
.B(n_227),
.C(n_226),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_583),
.A2(n_446),
.B(n_452),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_580),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_581),
.B(n_443),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_574),
.B(n_239),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_581),
.B(n_443),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_482),
.B(n_247),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_587),
.B(n_253),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_535),
.A2(n_219),
.B1(n_234),
.B2(n_237),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_587),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_507),
.A2(n_295),
.B1(n_243),
.B2(n_249),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_557),
.A2(n_250),
.B1(n_287),
.B2(n_298),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_590),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_491),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_541),
.B(n_297),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_480),
.A2(n_298),
.B1(n_287),
.B2(n_307),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_590),
.B(n_307),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_592),
.B(n_257),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_592),
.B(n_445),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_480),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_L g739 ( 
.A(n_561),
.B(n_442),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_595),
.B(n_445),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_598),
.B(n_445),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_596),
.B(n_262),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_527),
.A2(n_203),
.B1(n_445),
.B2(n_448),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_598),
.Y(n_744)
);

BUFx8_ASAP7_75t_L g745 ( 
.A(n_559),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_491),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_565),
.B(n_445),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_602),
.B(n_362),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_501),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_565),
.B(n_448),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_569),
.B(n_448),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_569),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_469),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_576),
.B(n_448),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_527),
.A2(n_203),
.B1(n_299),
.B2(n_292),
.Y(n_755)
);

NOR3xp33_ASAP7_75t_L g756 ( 
.A(n_614),
.B(n_566),
.C(n_561),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_609),
.B(n_576),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_647),
.B(n_558),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_611),
.A2(n_608),
.B(n_641),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_615),
.B(n_582),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_626),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_606),
.A2(n_582),
.B(n_594),
.C(n_593),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_635),
.A2(n_585),
.B(n_551),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_640),
.B(n_558),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_637),
.A2(n_617),
.B(n_662),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_629),
.B(n_518),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_629),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_606),
.B(n_290),
.C(n_263),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_643),
.A2(n_571),
.B1(n_575),
.B2(n_597),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_SL g770 ( 
.A1(n_707),
.A2(n_699),
.B(n_714),
.C(n_646),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_593),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_623),
.B(n_594),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_694),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_633),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_694),
.B(n_643),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_666),
.A2(n_585),
.B(n_521),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_618),
.A2(n_585),
.B(n_521),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_703),
.B(n_604),
.Y(n_778)
);

AOI21x1_ASAP7_75t_L g779 ( 
.A1(n_654),
.A2(n_605),
.B(n_604),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_629),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_636),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_665),
.B(n_527),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_627),
.A2(n_521),
.B(n_554),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_651),
.A2(n_521),
.B(n_554),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_642),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_645),
.Y(n_786)
);

NAND2x1p5_ASAP7_75t_L g787 ( 
.A(n_629),
.B(n_518),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_649),
.B(n_591),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_645),
.B(n_604),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_648),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_650),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_749),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_752),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_664),
.A2(n_605),
.B(n_493),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_708),
.A2(n_591),
.B1(n_518),
.B2(n_568),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_670),
.B(n_362),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_638),
.B(n_274),
.C(n_282),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_664),
.A2(n_563),
.B(n_551),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_676),
.A2(n_696),
.B(n_688),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_612),
.B(n_273),
.C(n_266),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_609),
.A2(n_527),
.B1(n_579),
.B2(n_568),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_742),
.B(n_264),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_673),
.B(n_527),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_638),
.A2(n_547),
.B(n_539),
.C(n_586),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_610),
.Y(n_805)
);

CKINVDCx8_ASAP7_75t_R g806 ( 
.A(n_705),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_677),
.B(n_547),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_749),
.B(n_468),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_674),
.A2(n_537),
.B(n_503),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_688),
.A2(n_563),
.B(n_551),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_678),
.A2(n_683),
.B1(n_691),
.B2(n_686),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_696),
.A2(n_493),
.B(n_563),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_697),
.B(n_468),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_704),
.A2(n_517),
.B1(n_468),
.B2(n_586),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_670),
.B(n_267),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_718),
.B(n_468),
.Y(n_816)
);

AOI33xp33_ASAP7_75t_L g817 ( 
.A1(n_616),
.A2(n_369),
.A3(n_363),
.B1(n_364),
.B2(n_366),
.B3(n_367),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_716),
.B(n_363),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_721),
.B(n_495),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_711),
.A2(n_712),
.B(n_720),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_728),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_731),
.B(n_495),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_659),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_712),
.A2(n_511),
.B(n_599),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_668),
.A2(n_579),
.B1(n_203),
.B2(n_506),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_675),
.A2(n_546),
.B(n_503),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_744),
.B(n_495),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_619),
.A2(n_546),
.B(n_523),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_749),
.B(n_495),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_632),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_624),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_693),
.A2(n_289),
.B(n_291),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_609),
.B(n_517),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_710),
.B(n_624),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_702),
.A2(n_511),
.B(n_599),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_682),
.A2(n_511),
.B(n_599),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_630),
.A2(n_528),
.B(n_523),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_709),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_607),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_634),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_690),
.B(n_275),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_619),
.A2(n_550),
.B(n_506),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_684),
.A2(n_497),
.B(n_599),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_609),
.B(n_517),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_693),
.A2(n_586),
.B(n_517),
.C(n_556),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_609),
.B(n_539),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_609),
.B(n_539),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_687),
.A2(n_511),
.B(n_497),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_723),
.B(n_364),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_723),
.B(n_276),
.C(n_310),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_692),
.A2(n_497),
.B(n_504),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_634),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_706),
.A2(n_497),
.B(n_504),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_668),
.A2(n_539),
.B1(n_586),
.B2(n_549),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_726),
.B(n_549),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_726),
.B(n_549),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_736),
.B(n_556),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_736),
.B(n_556),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_656),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_735),
.B(n_556),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_717),
.A2(n_532),
.B(n_504),
.Y(n_861)
);

BUFx4f_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_735),
.B(n_528),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_690),
.B(n_286),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_713),
.B(n_537),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_695),
.A2(n_550),
.B(n_560),
.C(n_544),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_713),
.B(n_538),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_722),
.A2(n_532),
.B(n_544),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_738),
.B(n_301),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_748),
.B(n_538),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_700),
.Y(n_871)
);

AOI33xp33_ASAP7_75t_L g872 ( 
.A1(n_616),
.A2(n_369),
.A3(n_366),
.B1(n_367),
.B2(n_442),
.B3(n_452),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_724),
.A2(n_532),
.B(n_560),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_679),
.A2(n_446),
.B(n_454),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_738),
.A2(n_451),
.B(n_452),
.C(n_454),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_622),
.A2(n_579),
.B(n_601),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_655),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_L g878 ( 
.A(n_695),
.B(n_308),
.C(n_454),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_737),
.A2(n_424),
.B(n_432),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_740),
.A2(n_424),
.B(n_432),
.Y(n_880)
);

BUFx2_ASAP7_75t_SL g881 ( 
.A(n_739),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_741),
.A2(n_432),
.B(n_446),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_628),
.B(n_579),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_644),
.B(n_579),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_671),
.B(n_579),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_671),
.A2(n_451),
.B(n_446),
.C(n_448),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_700),
.B(n_448),
.Y(n_887)
);

AND3x1_ASAP7_75t_L g888 ( 
.A(n_685),
.B(n_451),
.C(n_300),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_730),
.A2(n_448),
.B(n_432),
.C(n_300),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_681),
.B(n_3),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_639),
.B(n_709),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_622),
.B(n_579),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_747),
.A2(n_432),
.B(n_601),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_700),
.B(n_755),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_634),
.B(n_432),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_750),
.A2(n_432),
.B(n_601),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_657),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_733),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_700),
.B(n_601),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_660),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_620),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_753),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_625),
.Y(n_903)
);

BUFx8_ASAP7_75t_L g904 ( 
.A(n_634),
.Y(n_904)
);

OAI21xp33_ASAP7_75t_L g905 ( 
.A1(n_681),
.A2(n_6),
.B(n_7),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_613),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_680),
.A2(n_601),
.B(n_150),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_652),
.A2(n_755),
.B(n_727),
.C(n_658),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_661),
.B(n_9),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_701),
.B(n_9),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_631),
.A2(n_601),
.B(n_149),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_634),
.A2(n_601),
.B1(n_137),
.B2(n_134),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_653),
.B(n_10),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_733),
.A2(n_15),
.B(n_19),
.C(n_20),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_725),
.B(n_107),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_685),
.A2(n_20),
.B(n_27),
.C(n_32),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_667),
.Y(n_917)
);

BUFx12f_ASAP7_75t_L g918 ( 
.A(n_745),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_669),
.B(n_33),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_672),
.B(n_689),
.Y(n_920)
);

AO21x1_ASAP7_75t_L g921 ( 
.A1(n_751),
.A2(n_33),
.B(n_34),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_732),
.A2(n_133),
.B(n_131),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_773),
.B(n_831),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_764),
.B(n_831),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_R g925 ( 
.A(n_806),
.B(n_734),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_774),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_781),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_871),
.A2(n_754),
.B(n_700),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_786),
.B(n_734),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_775),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_786),
.B(n_815),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_805),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_839),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_760),
.A2(n_698),
.B1(n_663),
.B2(n_729),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_815),
.A2(n_719),
.B1(n_746),
.B2(n_700),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_906),
.B(n_35),
.Y(n_937)
);

OR2x2_ASAP7_75t_SL g938 ( 
.A(n_802),
.B(n_36),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_890),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_834),
.B(n_38),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_890),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_797),
.B(n_743),
.Y(n_942)
);

BUFx2_ASAP7_75t_SL g943 ( 
.A(n_788),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_871),
.A2(n_76),
.B(n_123),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_768),
.A2(n_128),
.B1(n_120),
.B2(n_116),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_796),
.B(n_46),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_849),
.B(n_47),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_780),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_758),
.B(n_805),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_902),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_768),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_878),
.A2(n_789),
.B(n_910),
.C(n_800),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_818),
.B(n_53),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_772),
.B(n_53),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_841),
.B(n_55),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_862),
.B(n_83),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_902),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_785),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_SL g959 ( 
.A(n_850),
.B(n_55),
.C(n_57),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_780),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_780),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_790),
.B(n_58),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_823),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_910),
.A2(n_61),
.B(n_88),
.C(n_93),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_850),
.B(n_101),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_918),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_790),
.B(n_105),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_905),
.B(n_869),
.C(n_832),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_SL g969 ( 
.A(n_869),
.B(n_864),
.C(n_841),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_859),
.B(n_891),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_789),
.A2(n_894),
.B1(n_885),
.B2(n_811),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_894),
.A2(n_799),
.B(n_762),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_778),
.B(n_791),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_759),
.A2(n_777),
.B(n_765),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_891),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_771),
.B(n_838),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_763),
.A2(n_776),
.B(n_887),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_878),
.B(n_756),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_794),
.A2(n_908),
.B(n_883),
.C(n_804),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_840),
.B(n_852),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_840),
.B(n_852),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_887),
.A2(n_833),
.B(n_847),
.Y(n_982)
);

AO21x1_ASAP7_75t_L g983 ( 
.A1(n_855),
.A2(n_858),
.B(n_857),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_821),
.A2(n_803),
.B(n_782),
.C(n_856),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_SL g985 ( 
.A1(n_907),
.A2(n_922),
.B(n_875),
.C(n_767),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_870),
.B(n_769),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_780),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_862),
.B(n_904),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_874),
.A2(n_837),
.B(n_783),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_L g990 ( 
.A(n_913),
.B(n_916),
.C(n_888),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_921),
.A2(n_825),
.B1(n_793),
.B2(n_917),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_767),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_844),
.A2(n_846),
.B(n_798),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_757),
.A2(n_779),
.B(n_784),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_757),
.A2(n_866),
.B(n_845),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_872),
.B(n_863),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_840),
.B(n_852),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_915),
.A2(n_881),
.B1(n_867),
.B2(n_865),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_840),
.B(n_852),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_877),
.B(n_897),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_915),
.B(n_825),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_859),
.B(n_792),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_900),
.B(n_817),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_901),
.A2(n_903),
.B1(n_860),
.B2(n_909),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_920),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_SL g1007 ( 
.A1(n_792),
.A2(n_876),
.B(n_809),
.C(n_826),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_L g1008 ( 
.A1(n_886),
.A2(n_889),
.B(n_835),
.C(n_814),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_810),
.A2(n_812),
.B(n_770),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_909),
.A2(n_919),
.B1(n_904),
.B2(n_807),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_898),
.A2(n_914),
.B(n_816),
.C(n_819),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_813),
.A2(n_827),
.B(n_822),
.C(n_854),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_795),
.B(n_884),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_766),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_892),
.A2(n_801),
.B(n_868),
.C(n_873),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_787),
.B(n_895),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_787),
.B(n_808),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_829),
.A2(n_824),
.B1(n_861),
.B2(n_836),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_829),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_828),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_911),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_842),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_899),
.B(n_843),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_SL g1024 ( 
.A1(n_848),
.A2(n_851),
.B(n_853),
.C(n_896),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_882),
.A2(n_912),
.B(n_893),
.C(n_880),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_899),
.B(n_879),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_761),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_780),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_773),
.B(n_615),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_773),
.B(n_615),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_764),
.B(n_615),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_764),
.B(n_615),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_775),
.A2(n_615),
.B1(n_773),
.B2(n_831),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_773),
.B(n_615),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_764),
.B(n_615),
.Y(n_1035)
);

NAND2x1_ASAP7_75t_L g1036 ( 
.A(n_780),
.B(n_767),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_806),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_890),
.A2(n_615),
.B1(n_905),
.B2(n_764),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_780),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_890),
.A2(n_615),
.B(n_815),
.C(n_606),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_780),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_871),
.A2(n_759),
.B(n_777),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_871),
.A2(n_759),
.B(n_777),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_780),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_775),
.A2(n_615),
.B1(n_773),
.B2(n_831),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_761),
.Y(n_1046)
);

AO21x1_ASAP7_75t_L g1047 ( 
.A1(n_890),
.A2(n_894),
.B(n_878),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_773),
.B(n_615),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_902),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_780),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_773),
.B(n_615),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_871),
.A2(n_759),
.B(n_777),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_806),
.B(n_649),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_890),
.A2(n_615),
.B(n_815),
.C(n_606),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_764),
.B(n_615),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_871),
.A2(n_759),
.B(n_777),
.Y(n_1056)
);

AOI22x1_ASAP7_75t_L g1057 ( 
.A1(n_799),
.A2(n_820),
.B1(n_834),
.B2(n_699),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_871),
.A2(n_759),
.B(n_777),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_932),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_933),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_960),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_933),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_925),
.B(n_1031),
.Y(n_1063)
);

AO31x2_ASAP7_75t_L g1064 ( 
.A1(n_1047),
.A2(n_983),
.A3(n_971),
.B(n_1056),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1035),
.B(n_1055),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_979),
.A2(n_986),
.B(n_984),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_993),
.A2(n_1009),
.B(n_928),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_950),
.Y(n_1071)
);

BUFx5_ASAP7_75t_L g1072 ( 
.A(n_1021),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1034),
.B(n_1048),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1052),
.A2(n_1058),
.B(n_982),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_1025),
.A2(n_1018),
.A3(n_1015),
.B(n_1023),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_958),
.Y(n_1076)
);

AO22x2_ASAP7_75t_L g1077 ( 
.A1(n_1002),
.A2(n_959),
.B1(n_990),
.B2(n_955),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1051),
.B(n_923),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_930),
.A2(n_972),
.B(n_985),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_975),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_1037),
.Y(n_1081)
);

AO22x1_ASAP7_75t_L g1082 ( 
.A1(n_937),
.A2(n_924),
.B1(n_940),
.B2(n_967),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_929),
.A2(n_1038),
.B1(n_973),
.B2(n_991),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_969),
.A2(n_1038),
.B(n_968),
.C(n_952),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_960),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_1026),
.A2(n_1033),
.A3(n_1045),
.B(n_1020),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1007),
.A2(n_1057),
.B(n_1012),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_995),
.A2(n_1008),
.B(n_1016),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_939),
.A2(n_941),
.B(n_951),
.C(n_937),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_940),
.B(n_1006),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_996),
.B(n_968),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_L g1092 ( 
.A(n_963),
.B(n_957),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_947),
.B(n_946),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_935),
.A2(n_1004),
.A3(n_953),
.B(n_944),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_964),
.B(n_998),
.C(n_965),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_954),
.A2(n_967),
.A3(n_1001),
.B(n_999),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1049),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1027),
.B(n_1046),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_942),
.A2(n_1011),
.B(n_936),
.C(n_991),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1053),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_925),
.B(n_1053),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_970),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1022),
.A2(n_1024),
.B(n_945),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_966),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_962),
.A2(n_934),
.A3(n_927),
.B(n_926),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_976),
.B(n_1003),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1005),
.A2(n_1017),
.B(n_997),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1010),
.A2(n_938),
.B1(n_981),
.B2(n_980),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1000),
.A2(n_981),
.B(n_980),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1014),
.B(n_943),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_1019),
.A2(n_1014),
.B(n_956),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1019),
.B(n_992),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1036),
.A2(n_948),
.B(n_1041),
.C(n_1028),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_988),
.A2(n_956),
.B1(n_992),
.B2(n_961),
.C(n_987),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_992),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_988),
.A2(n_1041),
.B(n_961),
.Y(n_1116)
);

AOI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_987),
.A2(n_1028),
.B1(n_960),
.B2(n_1039),
.C(n_1044),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_960),
.B(n_1039),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_1050),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1044),
.A2(n_974),
.B(n_1042),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1050),
.A2(n_974),
.B(n_1042),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1050),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_1040),
.B(n_1054),
.C(n_932),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_932),
.B(n_1031),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1040),
.B(n_1054),
.C(n_932),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_963),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_949),
.B(n_758),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_979),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_979),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_932),
.B(n_1031),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_970),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_1033),
.A2(n_1045),
.A3(n_971),
.B1(n_811),
.B2(n_1018),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_933),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_979),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_960),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_932),
.B(n_1031),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1141)
);

AOI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1013),
.A2(n_994),
.B(n_978),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_931),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_932),
.A2(n_615),
.B1(n_764),
.B2(n_1031),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1047),
.A2(n_983),
.A3(n_971),
.B(n_1042),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_932),
.B(n_834),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1053),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_932),
.A2(n_615),
.B1(n_1030),
.B2(n_1029),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_L g1150 ( 
.A(n_1040),
.B(n_1054),
.C(n_932),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_979),
.A2(n_972),
.B(n_995),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_992),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1154)
);

BUFx4_ASAP7_75t_SL g1155 ( 
.A(n_966),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_933),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1157)
);

AO32x2_ASAP7_75t_L g1158 ( 
.A1(n_1033),
.A2(n_1045),
.A3(n_971),
.B1(n_811),
.B2(n_1018),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_931),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1013),
.A2(n_994),
.B(n_978),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_932),
.B(n_1031),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_1053),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_931),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_960),
.B(n_1039),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_979),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_932),
.B(n_1031),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1040),
.B(n_1054),
.C(n_932),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_960),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_932),
.B(n_834),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_931),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_979),
.A2(n_972),
.B(n_995),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_974),
.A2(n_1043),
.B(n_1042),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_952),
.A2(n_1054),
.B(n_1040),
.C(n_1002),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_932),
.B(n_1031),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_989),
.A2(n_874),
.B(n_977),
.Y(n_1183)
);

INVx8_ASAP7_75t_L g1184 ( 
.A(n_1061),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1106),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1081),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1155),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1134),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1134),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1172),
.A2(n_1066),
.B1(n_1065),
.B2(n_1082),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1098),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1125),
.A2(n_1133),
.B1(n_1140),
.B2(n_1182),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1125),
.A2(n_1182),
.B1(n_1133),
.B2(n_1162),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1128),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1144),
.A2(n_1173),
.B1(n_1126),
.B2(n_1124),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_1104),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1060),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1176),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1062),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1156),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1140),
.A2(n_1162),
.B1(n_1157),
.B2(n_1168),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1076),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1124),
.A2(n_1126),
.B1(n_1173),
.B2(n_1150),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1063),
.A2(n_1078),
.B1(n_1149),
.B2(n_1073),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1129),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1150),
.A2(n_1069),
.B1(n_1073),
.B2(n_1078),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1077),
.A2(n_1095),
.B1(n_1149),
.B2(n_1130),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1089),
.A2(n_1077),
.B(n_1059),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1130),
.A2(n_1171),
.B1(n_1131),
.B2(n_1137),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1143),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1069),
.B(n_1090),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_1100),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1061),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1160),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1163),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1166),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_1080),
.Y(n_1217)
);

INVx6_ASAP7_75t_L g1218 ( 
.A(n_1061),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1061),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1146),
.B(n_1175),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1119),
.B(n_1174),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_SL g1222 ( 
.A(n_1102),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1095),
.A2(n_1171),
.B1(n_1131),
.B2(n_1137),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1093),
.B(n_1091),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_1148),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1083),
.A2(n_1067),
.B1(n_1151),
.B2(n_1177),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1085),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1083),
.A2(n_1067),
.B1(n_1151),
.B2(n_1177),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1103),
.A2(n_1108),
.B1(n_1101),
.B2(n_1079),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_1138),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1136),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_1071),
.B1(n_1110),
.B2(n_1097),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1153),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1115),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1099),
.A2(n_1092),
.B1(n_1108),
.B2(n_1107),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1103),
.A2(n_1107),
.B1(n_1087),
.B2(n_1111),
.Y(n_1236)
);

CKINVDCx11_ASAP7_75t_R g1237 ( 
.A(n_1138),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_1117),
.B1(n_1112),
.B2(n_1113),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1118),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1153),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1111),
.A2(n_1088),
.B1(n_1181),
.B2(n_1116),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1118),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1116),
.A2(n_1072),
.B1(n_1158),
.B2(n_1135),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1142),
.A2(n_1161),
.B1(n_1158),
.B2(n_1135),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1072),
.A2(n_1135),
.B1(n_1158),
.B2(n_1121),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1122),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1072),
.A2(n_1120),
.B1(n_1165),
.B2(n_1179),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1072),
.A2(n_1141),
.B1(n_1164),
.B2(n_1178),
.Y(n_1248)
);

BUFx8_ASAP7_75t_SL g1249 ( 
.A(n_1170),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1170),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1072),
.A2(n_1070),
.B1(n_1127),
.B2(n_1147),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1109),
.A2(n_1074),
.B1(n_1068),
.B2(n_1075),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1105),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1096),
.A2(n_1075),
.B1(n_1086),
.B2(n_1094),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1086),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1075),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1094),
.A2(n_1064),
.B1(n_1145),
.B2(n_1132),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1094),
.B(n_1064),
.Y(n_1258)
);

BUFx2_ASAP7_75t_SL g1259 ( 
.A(n_1145),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1145),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1123),
.A2(n_1139),
.B1(n_1152),
.B2(n_1154),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_SL g1262 ( 
.A(n_1159),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1167),
.A2(n_1169),
.B1(n_1180),
.B2(n_1183),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1061),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1098),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1125),
.A2(n_1140),
.B1(n_1162),
.B2(n_1133),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1125),
.A2(n_1140),
.B1(n_1162),
.B2(n_1133),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1129),
.B(n_758),
.Y(n_1269)
);

INVx6_ASAP7_75t_L g1270 ( 
.A(n_1061),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1106),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1061),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1172),
.A2(n_932),
.B1(n_1066),
.B2(n_1065),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

INVx8_ASAP7_75t_L g1279 ( 
.A(n_1061),
.Y(n_1279)
);

AOI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_1040),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1081),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1125),
.A2(n_1140),
.B1(n_1162),
.B2(n_1133),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1061),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1098),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1257),
.A2(n_1254),
.A3(n_1260),
.B(n_1255),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1253),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1223),
.B(n_1209),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1249),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1242),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1211),
.B(n_1224),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1209),
.A2(n_1236),
.B(n_1258),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1272),
.B(n_1275),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1239),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1256),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1256),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1280),
.A2(n_1208),
.B(n_1244),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1235),
.B(n_1259),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1261),
.A2(n_1263),
.B(n_1247),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1197),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1262),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1216),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1203),
.A2(n_1195),
.B(n_1207),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1203),
.B(n_1195),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1202),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1210),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1214),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1244),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1243),
.B(n_1226),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1221),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1236),
.A2(n_1245),
.B(n_1228),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1199),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1228),
.B(n_1220),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1193),
.B(n_1191),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1240),
.Y(n_1317)
);

BUFx8_ASAP7_75t_L g1318 ( 
.A(n_1186),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1265),
.Y(n_1319)
);

AOI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1238),
.A2(n_1232),
.B(n_1284),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1200),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1190),
.A2(n_1204),
.B1(n_1192),
.B2(n_1189),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1206),
.B(n_1229),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1231),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1206),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1273),
.B(n_1205),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1245),
.A2(n_1241),
.B(n_1248),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1184),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1229),
.B(n_1198),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1241),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1184),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1234),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1269),
.B(n_1185),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1267),
.A2(n_1271),
.B(n_1201),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1252),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1266),
.Y(n_1336)
);

INVx11_ASAP7_75t_L g1337 ( 
.A(n_1217),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1250),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1268),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

AO21x1_ASAP7_75t_L g1341 ( 
.A1(n_1282),
.A2(n_1201),
.B(n_1274),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1248),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1251),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1251),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1215),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1279),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1261),
.A2(n_1263),
.B(n_1247),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1213),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1218),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1187),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1219),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1233),
.B(n_1188),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1264),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1304),
.A2(n_1278),
.B1(n_1188),
.B2(n_1189),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1290),
.B(n_1316),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1338),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1345),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_R g1358 ( 
.A(n_1350),
.B(n_1227),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1300),
.A2(n_1283),
.B(n_1270),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_SL g1360 ( 
.A1(n_1304),
.A2(n_1334),
.B(n_1325),
.C(n_1353),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1326),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1316),
.B(n_1246),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1315),
.B(n_1194),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1289),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1333),
.B(n_1237),
.Y(n_1365)
);

NOR2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1288),
.B(n_1186),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1299),
.B(n_1281),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1312),
.B(n_1302),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1305),
.B(n_1278),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1305),
.B(n_1222),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1287),
.A2(n_1230),
.B(n_1283),
.C(n_1219),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1303),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1299),
.B(n_1219),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1306),
.B(n_1212),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1307),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1334),
.A2(n_1212),
.B1(n_1225),
.B2(n_1196),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1292),
.A2(n_1293),
.B1(n_1287),
.B2(n_1297),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1303),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1337),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1323),
.B(n_1320),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1310),
.A2(n_1325),
.B(n_1322),
.C(n_1336),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1310),
.A2(n_1336),
.B(n_1339),
.C(n_1340),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1301),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1320),
.A2(n_1339),
.B(n_1340),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1300),
.A2(n_1347),
.B(n_1330),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1314),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1329),
.B(n_1324),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1317),
.Y(n_1388)
);

AOI221xp5_ASAP7_75t_L g1389 ( 
.A1(n_1341),
.A2(n_1330),
.B1(n_1309),
.B2(n_1298),
.C(n_1321),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1329),
.B(n_1321),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1312),
.B(n_1302),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1341),
.B(n_1332),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1318),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1352),
.B(n_1319),
.Y(n_1394)
);

AOI221x1_ASAP7_75t_L g1395 ( 
.A1(n_1335),
.A2(n_1309),
.B1(n_1349),
.B2(n_1351),
.C(n_1348),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1311),
.B(n_1308),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1308),
.B(n_1291),
.Y(n_1397)
);

AND2x2_ASAP7_75t_SL g1398 ( 
.A(n_1313),
.B(n_1327),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1372),
.Y(n_1399)
);

INVx8_ASAP7_75t_L g1400 ( 
.A(n_1373),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1396),
.B(n_1298),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1398),
.B(n_1327),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1397),
.B(n_1285),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1396),
.B(n_1298),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_SL g1405 ( 
.A(n_1393),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1398),
.B(n_1397),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1359),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1359),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1385),
.B(n_1327),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1389),
.B(n_1298),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1327),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1385),
.B(n_1378),
.Y(n_1412)
);

INVx2_ASAP7_75t_R g1413 ( 
.A(n_1375),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1380),
.B(n_1342),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1392),
.B(n_1343),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1387),
.B(n_1285),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1392),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1390),
.B(n_1285),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1355),
.A2(n_1294),
.B1(n_1313),
.B2(n_1291),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1393),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1364),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1360),
.A2(n_1313),
.B1(n_1291),
.B2(n_1299),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1394),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1377),
.A2(n_1299),
.B1(n_1313),
.B2(n_1344),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1356),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1384),
.B(n_1291),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1425),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1403),
.B(n_1388),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1412),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1399),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1417),
.B(n_1394),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1403),
.B(n_1401),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1417),
.B(n_1414),
.Y(n_1433)
);

OAI31xp33_ASAP7_75t_L g1434 ( 
.A1(n_1410),
.A2(n_1381),
.A3(n_1360),
.B(n_1377),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1424),
.A2(n_1376),
.B1(n_1367),
.B2(n_1354),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1414),
.B(n_1382),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1424),
.A2(n_1381),
.B1(n_1376),
.B2(n_1369),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1410),
.A2(n_1362),
.B1(n_1370),
.B2(n_1371),
.C(n_1382),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1420),
.B(n_1361),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1415),
.B(n_1295),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1406),
.B(n_1368),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_1368),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1400),
.B(n_1367),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1412),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1395),
.C(n_1386),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1399),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_1391),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1415),
.B(n_1295),
.Y(n_1449)
);

AND2x2_ASAP7_75t_SL g1450 ( 
.A(n_1402),
.B(n_1286),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1399),
.Y(n_1451)
);

AND2x2_ASAP7_75t_SL g1452 ( 
.A(n_1426),
.B(n_1286),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1423),
.B(n_1404),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1423),
.B(n_1296),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1404),
.B(n_1285),
.Y(n_1457)
);

NOR3xp33_ASAP7_75t_L g1458 ( 
.A(n_1426),
.B(n_1383),
.C(n_1369),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1399),
.Y(n_1459)
);

AND3x1_ASAP7_75t_L g1460 ( 
.A(n_1405),
.B(n_1365),
.C(n_1371),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_SL g1461 ( 
.A(n_1419),
.B(n_1374),
.C(n_1363),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1443),
.B(n_1413),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1442),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1430),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1436),
.B(n_1421),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1433),
.B(n_1416),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1433),
.B(n_1416),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1447),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1443),
.B(n_1413),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1444),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1407),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1407),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1429),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1436),
.B(n_1416),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1407),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1442),
.B(n_1408),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1447),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1429),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1442),
.B(n_1408),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1429),
.B(n_1408),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1447),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1451),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1451),
.Y(n_1484)
);

OAI21xp33_ASAP7_75t_L g1485 ( 
.A1(n_1437),
.A2(n_1422),
.B(n_1411),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1418),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1451),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1440),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1453),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1459),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1409),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1459),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1432),
.B(n_1418),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1468),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1490),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1468),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1464),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_L g1501 ( 
.A(n_1485),
.B(n_1438),
.C(n_1446),
.Y(n_1501)
);

OAI32xp33_ASAP7_75t_L g1502 ( 
.A1(n_1485),
.A2(n_1446),
.A3(n_1457),
.B1(n_1438),
.B2(n_1432),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1464),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1465),
.B(n_1431),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1491),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1486),
.B(n_1434),
.C(n_1437),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1491),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1471),
.B(n_1448),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1469),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1465),
.B(n_1431),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1469),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1471),
.B(n_1450),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1475),
.B(n_1466),
.Y(n_1514)
);

NOR2x1p5_ASAP7_75t_L g1515 ( 
.A(n_1471),
.B(n_1420),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1471),
.B(n_1460),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1434),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1440),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1466),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1469),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1482),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1471),
.B(n_1448),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1467),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1489),
.A2(n_1461),
.B(n_1435),
.C(n_1452),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1439),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1467),
.B(n_1449),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1463),
.B(n_1448),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1482),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1473),
.B(n_1441),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1482),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1461),
.C(n_1422),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1463),
.B(n_1452),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1488),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1449),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1488),
.Y(n_1538)
);

AO21x1_ASAP7_75t_L g1539 ( 
.A1(n_1472),
.A2(n_1455),
.B(n_1428),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1463),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1500),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1501),
.B(n_1472),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1503),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1463),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1516),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1517),
.B(n_1452),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1515),
.Y(n_1547)
);

OAI32xp33_ASAP7_75t_L g1548 ( 
.A1(n_1501),
.A2(n_1457),
.A3(n_1470),
.B1(n_1462),
.B2(n_1472),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1498),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1509),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1497),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1516),
.B(n_1463),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1504),
.B(n_1481),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1473),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1499),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1510),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.B(n_1473),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1498),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1520),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1511),
.B(n_1481),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1505),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1476),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1476),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1521),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1494),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1524),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1476),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1474),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1571),
.A2(n_1532),
.B1(n_1524),
.B2(n_1460),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1557),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1551),
.B(n_1519),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1579)
);

AOI21xp33_ASAP7_75t_L g1580 ( 
.A1(n_1545),
.A2(n_1502),
.B(n_1519),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1288),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1542),
.A2(n_1546),
.B(n_1564),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1542),
.A2(n_1564),
.B1(n_1547),
.B2(n_1563),
.Y(n_1583)
);

AOI21xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1547),
.A2(n_1357),
.B(n_1379),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1563),
.B(n_1523),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1570),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1565),
.A2(n_1526),
.B1(n_1490),
.B2(n_1529),
.C(n_1534),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1539),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1477),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1548),
.A2(n_1357),
.B(n_1379),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1556),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1553),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1506),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1568),
.A2(n_1450),
.B1(n_1444),
.B2(n_1494),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1477),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1548),
.A2(n_1508),
.B(n_1528),
.C(n_1420),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1557),
.Y(n_1601)
);

OAI322xp33_ASAP7_75t_L g1602 ( 
.A1(n_1579),
.A2(n_1556),
.A3(n_1568),
.B1(n_1543),
.B2(n_1572),
.C1(n_1569),
.C2(n_1560),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1593),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1576),
.A2(n_1528),
.B(n_1560),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1543),
.C(n_1559),
.Y(n_1605)
);

AOI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1580),
.A2(n_1544),
.B(n_1540),
.C(n_1562),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1578),
.A2(n_1562),
.B(n_1554),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1581),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1577),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1569),
.C(n_1561),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1594),
.A2(n_1450),
.B1(n_1540),
.B2(n_1544),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1596),
.A2(n_1570),
.B1(n_1566),
.B2(n_1567),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1600),
.A2(n_1554),
.B(n_1561),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1601),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1598),
.A2(n_1570),
.B1(n_1566),
.B2(n_1567),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1591),
.A2(n_1405),
.B1(n_1288),
.B2(n_1420),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1589),
.A2(n_1570),
.B1(n_1559),
.B2(n_1549),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1616),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1603),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1607),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1609),
.B(n_1586),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1627)
);

OAI31xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1611),
.A2(n_1608),
.A3(n_1605),
.B(n_1621),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1587),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1610),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1629),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_L g1634 ( 
.A(n_1626),
.B(n_1612),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1630),
.B(n_1602),
.Y(n_1635)
);

OAI21xp33_ASAP7_75t_L g1636 ( 
.A1(n_1628),
.A2(n_1613),
.B(n_1618),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1622),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1624),
.Y(n_1639)
);

OAI211xp5_ASAP7_75t_L g1640 ( 
.A1(n_1627),
.A2(n_1612),
.B(n_1614),
.C(n_1623),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1627),
.B(n_1625),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1632),
.A2(n_1620),
.B(n_1592),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1635),
.A2(n_1615),
.B(n_1590),
.Y(n_1644)
);

XNOR2xp5_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1366),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1635),
.A2(n_1585),
.B1(n_1599),
.B2(n_1601),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1633),
.A2(n_1599),
.B1(n_1559),
.B2(n_1574),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1640),
.A2(n_1572),
.B(n_1559),
.Y(n_1648)
);

AOI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1637),
.A2(n_1536),
.B(n_1533),
.Y(n_1649)
);

NAND2x1_ASAP7_75t_L g1650 ( 
.A(n_1647),
.B(n_1643),
.Y(n_1650)
);

AOI21xp33_ASAP7_75t_L g1651 ( 
.A1(n_1645),
.A2(n_1636),
.B(n_1634),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1646),
.A2(n_1641),
.B1(n_1638),
.B2(n_1574),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1648),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1644),
.A2(n_1642),
.B(n_1649),
.C(n_1549),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1644),
.A2(n_1575),
.B(n_1555),
.C(n_1573),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1653),
.B(n_1573),
.Y(n_1656)
);

NAND4xp75_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1318),
.C(n_1337),
.D(n_1558),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1650),
.A2(n_1558),
.B1(n_1575),
.B2(n_1538),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1654),
.B(n_1477),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1652),
.A2(n_1470),
.B(n_1462),
.Y(n_1660)
);

NAND4xp75_ASAP7_75t_L g1661 ( 
.A(n_1659),
.B(n_1655),
.C(n_1318),
.D(n_1358),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1657),
.B(n_1318),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1656),
.A2(n_1480),
.B1(n_1462),
.B2(n_1470),
.Y(n_1663)
);

AND3x4_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1658),
.C(n_1358),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1664),
.Y(n_1665)
);

XNOR2xp5_ASAP7_75t_L g1666 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1665),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1667),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1666),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1668),
.A2(n_1660),
.B1(n_1663),
.B2(n_1427),
.Y(n_1670)
);

OA22x2_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1474),
.B1(n_1479),
.B2(n_1480),
.Y(n_1671)
);

OAI322xp33_ASAP7_75t_L g1672 ( 
.A1(n_1670),
.A2(n_1495),
.A3(n_1478),
.B1(n_1483),
.B2(n_1484),
.C1(n_1493),
.C2(n_1479),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1672),
.B(n_1671),
.Y(n_1673)
);

XNOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1673),
.B(n_1346),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1495),
.B1(n_1346),
.B2(n_1427),
.C(n_1493),
.Y(n_1675)
);

AOI211xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1331),
.B(n_1328),
.C(n_1346),
.Y(n_1676)
);


endmodule