module real_aes_8662_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g441 ( .A(n_0), .Y(n_441) );
INVx1_ASAP7_75t_L g533 ( .A(n_1), .Y(n_533) );
INVx1_ASAP7_75t_L g151 ( .A(n_2), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_3), .A2(n_39), .B1(n_176), .B2(n_479), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g183 ( .A1(n_4), .A2(n_167), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_5), .B(n_165), .Y(n_545) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_7), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_8), .B(n_40), .Y(n_442) );
INVx1_ASAP7_75t_L g189 ( .A(n_9), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_10), .B(n_246), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_11), .A2(n_102), .B1(n_114), .B2(n_741), .Y(n_101) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_13), .B(n_157), .Y(n_488) );
INVx1_ASAP7_75t_L g260 ( .A(n_14), .Y(n_260) );
INVx1_ASAP7_75t_L g527 ( .A(n_15), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_16), .B(n_132), .Y(n_516) );
AO32x2_ASAP7_75t_L g500 ( .A1(n_17), .A2(n_131), .A3(n_165), .B1(n_481), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_18), .B(n_176), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_19), .B(n_172), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_20), .B(n_132), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_21), .A2(n_50), .B1(n_176), .B2(n_479), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_22), .B(n_167), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_23), .A2(n_97), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_23), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_24), .A2(n_75), .B1(n_157), .B2(n_176), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_25), .B(n_176), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_26), .B(n_179), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_27), .A2(n_258), .B(n_259), .C(n_261), .Y(n_257) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_28), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_29), .B(n_162), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_30), .B(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_31), .A2(n_87), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_31), .Y(n_122) );
INVx1_ASAP7_75t_L g204 ( .A(n_32), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_33), .B(n_162), .Y(n_472) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_34), .A2(n_447), .B1(n_731), .B2(n_732), .C1(n_735), .C2(n_737), .Y(n_446) );
INVx2_ASAP7_75t_L g142 ( .A(n_35), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_36), .B(n_176), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_37), .B(n_162), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_38), .A2(n_144), .B(n_147), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_40), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g202 ( .A(n_41), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_42), .B(n_155), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_43), .B(n_176), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_44), .A2(n_85), .B1(n_224), .B2(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_45), .B(n_176), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_46), .B(n_176), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_47), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_48), .B(n_532), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_49), .B(n_167), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_51), .A2(n_60), .B1(n_157), .B2(n_176), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_52), .A2(n_147), .B1(n_157), .B2(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_53), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_54), .B(n_176), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_55), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_56), .B(n_176), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_57), .A2(n_175), .B(n_187), .C(n_188), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_58), .Y(n_237) );
INVx1_ASAP7_75t_L g185 ( .A(n_59), .Y(n_185) );
INVx1_ASAP7_75t_L g145 ( .A(n_61), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_62), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_63), .B(n_176), .Y(n_534) );
INVx1_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
AO32x2_ASAP7_75t_L g476 ( .A1(n_66), .A2(n_165), .A3(n_240), .B1(n_477), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g552 ( .A(n_67), .Y(n_552) );
INVx1_ASAP7_75t_L g467 ( .A(n_68), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_69), .A2(n_172), .B(n_173), .C(n_175), .Y(n_171) );
INVxp67_ASAP7_75t_L g174 ( .A(n_70), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_71), .B(n_157), .Y(n_468) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_73), .Y(n_207) );
INVx1_ASAP7_75t_L g230 ( .A(n_74), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_76), .A2(n_144), .B(n_147), .C(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_77), .B(n_479), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_78), .B(n_157), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_79), .B(n_152), .Y(n_220) );
INVx2_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_81), .B(n_172), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_82), .B(n_157), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_83), .A2(n_144), .B(n_147), .C(n_150), .Y(n_146) );
INVx2_ASAP7_75t_L g110 ( .A(n_84), .Y(n_110) );
OR2x2_ASAP7_75t_L g438 ( .A(n_84), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g450 ( .A(n_84), .B(n_440), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_86), .A2(n_100), .B1(n_157), .B2(n_158), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_87), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_88), .B(n_162), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_89), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_90), .A2(n_144), .B(n_147), .C(n_243), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_91), .Y(n_250) );
INVx1_ASAP7_75t_L g170 ( .A(n_92), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_93), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_94), .B(n_152), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_95), .B(n_157), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_96), .B(n_165), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_97), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_99), .A2(n_167), .B(n_168), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g741 ( .A(n_104), .Y(n_741) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g454 ( .A(n_110), .B(n_440), .Y(n_454) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_110), .B(n_439), .Y(n_739) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_445), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g740 ( .A(n_116), .Y(n_740) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_436), .B(n_443), .Y(n_119) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx1_ASAP7_75t_L g451 ( .A(n_124), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_124), .A2(n_452), .B1(n_456), .B2(n_736), .Y(n_735) );
NAND2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_352), .Y(n_124) );
NOR5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_275), .C(n_307), .D(n_322), .E(n_339), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_191), .B(n_212), .C(n_263), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_163), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_128), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_128), .B(n_327), .Y(n_390) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_129), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_129), .B(n_209), .Y(n_276) );
AND2x2_ASAP7_75t_L g317 ( .A(n_129), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_129), .B(n_286), .Y(n_321) );
OR2x2_ASAP7_75t_L g358 ( .A(n_129), .B(n_197), .Y(n_358) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g196 ( .A(n_130), .B(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g266 ( .A(n_130), .Y(n_266) );
OR2x2_ASAP7_75t_L g429 ( .A(n_130), .B(n_269), .Y(n_429) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_137), .B(n_159), .Y(n_130) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_131), .A2(n_198), .B(n_206), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_131), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_133), .B(n_134), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_146), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_139), .A2(n_177), .B1(n_199), .B2(n_205), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_139), .A2(n_230), .B(n_231), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
AND2x4_ASAP7_75t_L g167 ( .A(n_140), .B(n_144), .Y(n_167) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g532 ( .A(n_141), .Y(n_532) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx3_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_143), .Y(n_155) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx4_ASAP7_75t_SL g177 ( .A(n_144), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_144), .A2(n_466), .B(n_469), .Y(n_465) );
BUFx3_ASAP7_75t_L g481 ( .A(n_144), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_144), .A2(n_486), .B(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_144), .A2(n_526), .B(n_530), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_144), .A2(n_539), .B(n_542), .Y(n_538) );
INVx5_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
BUFx3_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
INVx1_ASAP7_75t_L g479 ( .A(n_148), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_154), .C(n_156), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_SL g466 ( .A1(n_152), .A2(n_175), .B(n_467), .C(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g503 ( .A(n_152), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_152), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_152), .A2(n_549), .B(n_550), .Y(n_548) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_153), .B(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_153), .B(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g477 ( .A1(n_153), .A2(n_155), .B1(n_478), .B2(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx4_ASAP7_75t_L g246 ( .A(n_155), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_155), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_155), .A2(n_503), .B1(n_519), .B2(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_156), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_161), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_161), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_162), .A2(n_253), .B(n_262), .Y(n_252) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_162), .A2(n_465), .B(n_472), .Y(n_464) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_162), .A2(n_485), .B(n_493), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_163), .A2(n_332), .B1(n_333), .B2(n_336), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_163), .B(n_266), .Y(n_415) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_181), .Y(n_163) );
AND2x2_ASAP7_75t_L g211 ( .A(n_164), .B(n_197), .Y(n_211) );
AND2x2_ASAP7_75t_L g268 ( .A(n_164), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g273 ( .A(n_164), .Y(n_273) );
INVx3_ASAP7_75t_L g286 ( .A(n_164), .Y(n_286) );
OR2x2_ASAP7_75t_L g306 ( .A(n_164), .B(n_269), .Y(n_306) );
AND2x2_ASAP7_75t_L g325 ( .A(n_164), .B(n_182), .Y(n_325) );
BUFx2_ASAP7_75t_L g357 ( .A(n_164), .Y(n_357) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_178), .Y(n_164) );
INVx4_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_165), .A2(n_538), .B(n_545), .Y(n_537) );
BUFx2_ASAP7_75t_L g254 ( .A(n_167), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_177), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_169), .A2(n_177), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_169), .A2(n_177), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g489 ( .A(n_172), .Y(n_489) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_176), .Y(n_247) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_179), .A2(n_183), .B(n_190), .Y(n_182) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_180), .B(n_227), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_180), .B(n_481), .C(n_518), .Y(n_517) );
AO21x1_ASAP7_75t_L g607 ( .A1(n_180), .A2(n_518), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g272 ( .A(n_181), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
BUFx2_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
INVx2_ASAP7_75t_L g210 ( .A(n_182), .Y(n_210) );
OR2x2_ASAP7_75t_L g288 ( .A(n_182), .B(n_269), .Y(n_288) );
AND2x2_ASAP7_75t_L g318 ( .A(n_182), .B(n_197), .Y(n_318) );
AND2x2_ASAP7_75t_L g335 ( .A(n_182), .B(n_266), .Y(n_335) );
AND2x2_ASAP7_75t_L g375 ( .A(n_182), .B(n_286), .Y(n_375) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_182), .B(n_211), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_187), .A2(n_491), .B(n_492), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g551 ( .A1(n_187), .A2(n_531), .B(n_552), .C(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp33_ASAP7_75t_SL g192 ( .A(n_193), .B(n_208), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_194), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_195), .A2(n_211), .B(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_195), .B(n_197), .Y(n_405) );
AND2x2_ASAP7_75t_L g341 ( .A(n_196), .B(n_342), .Y(n_341) );
INVx3_ASAP7_75t_L g269 ( .A(n_197), .Y(n_269) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_197), .Y(n_367) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_200) );
INVx2_ASAP7_75t_L g203 ( .A(n_201), .Y(n_203) );
INVx4_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_208), .B(n_266), .Y(n_434) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_209), .A2(n_377), .B1(n_378), .B2(n_383), .Y(n_376) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AND2x2_ASAP7_75t_L g267 ( .A(n_210), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g342 ( .A(n_210), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_211), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g396 ( .A(n_211), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_238), .Y(n_213) );
INVx4_ASAP7_75t_L g282 ( .A(n_214), .Y(n_282) );
AND2x2_ASAP7_75t_L g360 ( .A(n_214), .B(n_327), .Y(n_360) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
INVx3_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_215), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_215), .Y(n_297) );
INVx2_ASAP7_75t_L g311 ( .A(n_215), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_215), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g368 ( .A(n_215), .B(n_363), .Y(n_368) );
AND2x2_ASAP7_75t_L g433 ( .A(n_215), .B(n_403), .Y(n_433) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_218), .B(n_225), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_222), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
INVx1_ASAP7_75t_L g235 ( .A(n_225), .Y(n_235) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_225), .A2(n_525), .B(n_535), .Y(n_524) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_225), .A2(n_547), .B(n_554), .Y(n_546) );
AND2x2_ASAP7_75t_L g274 ( .A(n_228), .B(n_252), .Y(n_274) );
INVx2_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_235), .B(n_236), .Y(n_228) );
INVx1_ASAP7_75t_L g299 ( .A(n_238), .Y(n_299) );
AND2x2_ASAP7_75t_L g345 ( .A(n_238), .B(n_293), .Y(n_345) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_251), .Y(n_238) );
INVx2_ASAP7_75t_L g284 ( .A(n_239), .Y(n_284) );
INVx1_ASAP7_75t_L g292 ( .A(n_239), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_239), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_239), .B(n_294), .Y(n_348) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_249), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_248), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_247), .Y(n_243) );
AND2x2_ASAP7_75t_L g327 ( .A(n_251), .B(n_284), .Y(n_327) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
AND2x2_ASAP7_75t_L g363 ( .A(n_252), .B(n_294), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_258), .B(n_260), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_258), .A2(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g529 ( .A(n_258), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_270), .B(n_274), .Y(n_263) );
INVx1_ASAP7_75t_SL g308 ( .A(n_264), .Y(n_308) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_265), .B(n_272), .Y(n_365) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g314 ( .A(n_266), .B(n_269), .Y(n_314) );
AND2x2_ASAP7_75t_L g343 ( .A(n_266), .B(n_287), .Y(n_343) );
OR2x2_ASAP7_75t_L g346 ( .A(n_266), .B(n_306), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_267), .A2(n_359), .B1(n_411), .B2(n_412), .C1(n_414), .C2(n_416), .Y(n_410) );
BUFx2_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_314), .Y(n_313) );
INVx3_ASAP7_75t_SL g330 ( .A(n_272), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_272), .B(n_324), .Y(n_384) );
AND2x2_ASAP7_75t_L g319 ( .A(n_274), .B(n_279), .Y(n_319) );
INVx1_ASAP7_75t_L g338 ( .A(n_274), .Y(n_338) );
OAI221xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_277), .B1(n_281), .B2(n_285), .C(n_289), .Y(n_275) );
OR2x2_ASAP7_75t_L g347 ( .A(n_277), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g332 ( .A(n_279), .B(n_302), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_279), .B(n_292), .Y(n_372) );
AND2x2_ASAP7_75t_L g377 ( .A(n_279), .B(n_327), .Y(n_377) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_279), .Y(n_387) );
NAND2x1_ASAP7_75t_SL g398 ( .A(n_279), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g283 ( .A(n_280), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_280), .B(n_298), .Y(n_329) );
INVx1_ASAP7_75t_L g395 ( .A(n_280), .Y(n_395) );
INVx1_ASAP7_75t_L g370 ( .A(n_281), .Y(n_370) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g382 ( .A(n_282), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_282), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g399 ( .A(n_283), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_283), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g302 ( .A(n_284), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_284), .B(n_294), .Y(n_315) );
INVx1_ASAP7_75t_L g381 ( .A(n_284), .Y(n_381) );
INVx1_ASAP7_75t_L g402 ( .A(n_285), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_295), .B(n_304), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g435 ( .A(n_291), .B(n_368), .Y(n_435) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g403 ( .A(n_292), .B(n_363), .Y(n_403) );
AOI32xp33_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_299), .A3(n_317), .B1(n_319), .B2(n_320), .Y(n_316) );
AOI322xp5_ASAP7_75t_L g418 ( .A1(n_293), .A2(n_325), .A3(n_408), .B1(n_419), .B2(n_420), .C1(n_421), .C2(n_423), .Y(n_418) );
INVx2_ASAP7_75t_L g298 ( .A(n_294), .Y(n_298) );
INVx1_ASAP7_75t_L g408 ( .A(n_294), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_300), .B2(n_301), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_296), .B(n_302), .Y(n_351) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_297), .B(n_363), .Y(n_413) );
INVx1_ASAP7_75t_L g300 ( .A(n_298), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_298), .B(n_327), .Y(n_417) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_306), .B(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_309), .B1(n_312), .B2(n_315), .C(n_316), .Y(n_307) );
OR2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g337 ( .A(n_309), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g362 ( .A(n_310), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g366 ( .A(n_320), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B1(n_328), .B2(n_330), .C(n_331), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_324), .A2(n_355), .B1(n_359), .B2(n_360), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_325), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_325), .Y(n_430) );
INVx1_ASAP7_75t_L g424 ( .A(n_327), .Y(n_424) );
INVx1_ASAP7_75t_SL g359 ( .A(n_328), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_330), .B(n_358), .Y(n_420) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_335), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g401 ( .A(n_335), .Y(n_401) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
OAI221xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_344), .B1(n_346), .B2(n_347), .C(n_349), .Y(n_339) );
NOR2xp33_ASAP7_75t_SL g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_341), .A2(n_359), .B1(n_405), .B2(n_406), .Y(n_404) );
CKINVDCx14_ASAP7_75t_R g344 ( .A(n_345), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g423 ( .A1(n_346), .A2(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_SL g352 ( .A(n_353), .B(n_385), .C(n_409), .Y(n_352) );
NAND4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_361), .C(n_369), .D(n_376), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
INVx3_ASAP7_75t_SL g426 ( .A(n_358), .Y(n_426) );
OR2x2_ASAP7_75t_L g431 ( .A(n_358), .B(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_366), .B2(n_368), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_363), .B(n_381), .Y(n_422) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B(n_373), .Y(n_369) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_391), .C(n_404), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_396), .B1(n_397), .B2(n_400), .C1(n_402), .C2(n_403), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND4xp25_ASAP7_75t_SL g428 ( .A(n_401), .B(n_429), .C(n_430), .D(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND3xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_418), .C(n_427), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_433), .B1(n_434), .B2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g444 ( .A(n_438), .Y(n_444) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_443), .A2(n_446), .B(n_740), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_452), .B2(n_455), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g736 ( .A(n_449), .Y(n_736) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_652), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_601), .C(n_643), .Y(n_457) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_510), .B(n_555), .C(n_577), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_473), .B(n_494), .C(n_505), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_461), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g664 ( .A(n_461), .B(n_581), .Y(n_664) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g566 ( .A(n_462), .B(n_497), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_462), .B(n_484), .Y(n_683) );
INVx1_ASAP7_75t_L g701 ( .A(n_462), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_462), .B(n_598), .Y(n_710) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g593 ( .A(n_463), .B(n_484), .Y(n_593) );
AND2x2_ASAP7_75t_L g651 ( .A(n_463), .B(n_598), .Y(n_651) );
INVx1_ASAP7_75t_L g695 ( .A(n_463), .Y(n_695) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g572 ( .A(n_464), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g580 ( .A(n_464), .Y(n_580) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_464), .Y(n_620) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .Y(n_474) );
AND2x2_ASAP7_75t_L g559 ( .A(n_475), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g592 ( .A(n_475), .Y(n_592) );
OR2x2_ASAP7_75t_L g718 ( .A(n_475), .B(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_475), .B(n_484), .Y(n_722) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g497 ( .A(n_476), .Y(n_497) );
INVx1_ASAP7_75t_L g508 ( .A(n_476), .Y(n_508) );
AND2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_499), .Y(n_581) );
AND2x2_ASAP7_75t_L g621 ( .A(n_476), .B(n_500), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_481), .A2(n_548), .B(n_551), .Y(n_547) );
INVxp67_ASAP7_75t_L g663 ( .A(n_482), .Y(n_663) );
AND2x4_ASAP7_75t_L g688 ( .A(n_482), .B(n_581), .Y(n_688) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_483), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g498 ( .A(n_484), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g567 ( .A(n_484), .B(n_500), .Y(n_567) );
INVx1_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
INVx2_ASAP7_75t_L g599 ( .A(n_484), .Y(n_599) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_616), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_495), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
AND2x2_ASAP7_75t_L g678 ( .A(n_497), .B(n_499), .Y(n_678) );
AND2x2_ASAP7_75t_L g595 ( .A(n_498), .B(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g694 ( .A(n_498), .B(n_695), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_499), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g719 ( .A(n_499), .B(n_580), .Y(n_719) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g509 ( .A(n_500), .Y(n_509) );
AND2x2_ASAP7_75t_L g598 ( .A(n_500), .B(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_503), .A2(n_531), .B(n_533), .C(n_534), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_503), .A2(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x2_ASAP7_75t_L g644 ( .A(n_507), .B(n_579), .Y(n_644) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_508), .B(n_580), .Y(n_629) );
INVx2_ASAP7_75t_L g628 ( .A(n_509), .Y(n_628) );
OAI222xp33_ASAP7_75t_L g632 ( .A1(n_509), .A2(n_572), .B1(n_633), .B2(n_635), .C1(n_636), .C2(n_639), .Y(n_632) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g557 ( .A(n_514), .Y(n_557) );
OR2x2_ASAP7_75t_L g668 ( .A(n_514), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_515), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g647 ( .A(n_515), .B(n_561), .Y(n_647) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g608 ( .A(n_516), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_521), .A2(n_611), .B1(n_650), .B2(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_536), .Y(n_521) );
INVx3_ASAP7_75t_L g583 ( .A(n_522), .Y(n_583) );
OR2x2_ASAP7_75t_L g716 ( .A(n_522), .B(n_592), .Y(n_716) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g605 ( .A(n_523), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g613 ( .A(n_523), .B(n_561), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_523), .B(n_537), .Y(n_669) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_524), .B(n_537), .Y(n_564) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_587), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_524), .B(n_546), .Y(n_680) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_536), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_557), .Y(n_596) );
AND2x2_ASAP7_75t_L g600 ( .A(n_536), .B(n_590), .Y(n_600) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_546), .Y(n_536) );
INVx3_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g721 ( .A(n_537), .B(n_704), .Y(n_721) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_546), .Y(n_575) );
INVx2_ASAP7_75t_L g587 ( .A(n_546), .Y(n_587) );
AND2x2_ASAP7_75t_L g631 ( .A(n_546), .B(n_607), .Y(n_631) );
INVx1_ASAP7_75t_L g674 ( .A(n_546), .Y(n_674) );
OR2x2_ASAP7_75t_L g705 ( .A(n_546), .B(n_607), .Y(n_705) );
AND2x2_ASAP7_75t_L g725 ( .A(n_546), .B(n_561), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g563 ( .A(n_557), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_557), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g682 ( .A(n_559), .Y(n_682) );
INVx2_ASAP7_75t_SL g576 ( .A(n_560), .Y(n_576) );
AND2x2_ASAP7_75t_L g696 ( .A(n_560), .B(n_590), .Y(n_696) );
INVx2_ASAP7_75t_L g642 ( .A(n_561), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_568), .B2(n_574), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_564), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g730 ( .A(n_564), .Y(n_730) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g655 ( .A(n_566), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_566), .B(n_598), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_567), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g671 ( .A(n_567), .B(n_620), .Y(n_671) );
INVx2_ASAP7_75t_L g727 ( .A(n_567), .Y(n_727) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g597 ( .A(n_570), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_570), .B(n_615), .Y(n_648) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_572), .B(n_592), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g709 ( .A(n_575), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_576), .A2(n_660), .B(n_662), .C(n_665), .Y(n_659) );
OR2x2_ASAP7_75t_L g686 ( .A(n_576), .B(n_590), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_582), .B1(n_584), .B2(n_591), .C(n_594), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_579), .B(n_628), .Y(n_635) );
AND2x2_ASAP7_75t_L g677 ( .A(n_579), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
INVx1_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_583), .B(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g691 ( .A(n_583), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_583), .B(n_631), .Y(n_707) );
INVx2_ASAP7_75t_L g693 ( .A(n_584), .Y(n_693) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g634 ( .A(n_586), .B(n_605), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_586), .A2(n_602), .B(n_644), .C(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g612 ( .A(n_587), .B(n_607), .Y(n_612) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_591), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g660 ( .A(n_592), .B(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_600), .Y(n_594) );
INVx1_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
INVx1_ASAP7_75t_L g661 ( .A(n_598), .Y(n_661) );
INVx1_ASAP7_75t_L g712 ( .A(n_600), .Y(n_712) );
AOI211xp5_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_605), .B(n_609), .C(n_632), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g624 ( .A(n_604), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g675 ( .A(n_605), .Y(n_675) );
AND2x2_ASAP7_75t_L g724 ( .A(n_605), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_614), .B(n_622), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g638 ( .A(n_612), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_612), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g630 ( .A(n_613), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g706 ( .A(n_613), .Y(n_706) );
OAI32xp33_ASAP7_75t_L g717 ( .A1(n_613), .A2(n_665), .A3(n_672), .B1(n_713), .B2(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_618), .Y(n_614) );
INVx1_ASAP7_75t_SL g685 ( .A(n_615), .Y(n_685) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g625 ( .A(n_621), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_630), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_624), .A2(n_672), .B1(n_698), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_628), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g658 ( .A(n_642), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B(n_649), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_651), .A2(n_693), .B1(n_694), .B2(n_696), .C(n_697), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g652 ( .A(n_653), .B(n_676), .C(n_692), .D(n_702), .E(n_720), .Y(n_652) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_659), .C(n_666), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g723 ( .A(n_660), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_670), .B2(n_672), .Y(n_666) );
INVx1_ASAP7_75t_SL g699 ( .A(n_669), .Y(n_699) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_672), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_681) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g684 ( .A(n_674), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_674), .B(n_699), .Y(n_698) );
AOI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_679), .B(n_681), .C(n_689), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_685), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g728 ( .A(n_695), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_710), .B1(n_711), .B2(n_715), .C(n_717), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_706), .B(n_707), .C(n_708), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g729 ( .A(n_705), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_720) );
AOI21xp33_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_728), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule