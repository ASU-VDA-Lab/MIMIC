module fake_jpeg_29478_n_53 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_21),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_7),
.B(n_16),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_8),
.B(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_23),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_22),
.B1(n_15),
.B2(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_11),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_1),
.C(n_2),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_33),
.C(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.C(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_40),
.B2(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_44),
.Y(n_50)
);

AOI321xp33_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_46),
.A3(n_48),
.B1(n_49),
.B2(n_6),
.C(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_4),
.B(n_5),
.Y(n_53)
);


endmodule