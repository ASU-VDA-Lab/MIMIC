module real_jpeg_19406_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_244;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_0),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_26),
.B1(n_60),
.B2(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_58),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_0),
.A2(n_10),
.B(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_0),
.B(n_126),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_0),
.A2(n_60),
.B(n_76),
.C(n_212),
.Y(n_211)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_3),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_3),
.B(n_176),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_5),
.A2(n_34),
.B1(n_60),
.B2(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_34),
.B1(n_55),
.B2(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_70),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_70),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_70),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_37),
.B(n_40),
.C(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_10),
.B(n_40),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_11),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_137),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_135),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_107),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_15),
.B(n_107),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_84),
.B2(n_85),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_21),
.B(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_22),
.B(n_30),
.Y(n_166)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_23),
.A2(n_31),
.B(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_24),
.B(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_26),
.A2(n_38),
.B(n_41),
.C(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_26),
.B(n_36),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_26),
.B(n_28),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_26),
.A2(n_40),
.B(n_77),
.Y(n_212)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_28),
.A2(n_29),
.B(n_95),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_30),
.B(n_176),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_31),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B(n_45),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_36),
.A2(n_89),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_37),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_37),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_37),
.B(n_99),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_39),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_41),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_45),
.B(n_183),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_47),
.B(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_71),
.B2(n_83),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_63),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_54),
.B(n_65),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_59),
.B(n_66),
.C(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_66),
.Y(n_67)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_69),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_75),
.B(n_76),
.C(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_62),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_61),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_73),
.B(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_74),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_81),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_78),
.B(n_150),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_80),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_86),
.A2(n_87),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_87),
.B(n_211),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_90),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.C(n_103),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_96),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_98),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_108),
.B(n_111),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_112),
.A2(n_113),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_123),
.C(n_131),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_115),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_124),
.B1(n_131),
.B2(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_244),
.C(n_249),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_156),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_156),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_153),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_141),
.B(n_142),
.C(n_153),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_148),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_157),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_162),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_163),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_175),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_243),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_237),
.B(n_242),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_222),
.B(n_236),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_207),
.B(n_221),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_196),
.B(n_206),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_185),
.B(n_195),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2x1_ASAP7_75t_R g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_215),
.B2(n_220),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_231),
.C(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule