module fake_aes_10901_n_41 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41, n_35);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
output n_35;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_2), .B(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_5), .B(n_7), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_16), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_13), .B(n_0), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_18), .B1(n_15), .B2(n_17), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_17), .B(n_18), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_23), .Y(n_29) );
AOI31xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_22), .A3(n_23), .B(n_15), .Y(n_30) );
NAND4xp25_ASAP7_75t_L g31 ( .A(n_28), .B(n_20), .C(n_15), .D(n_12), .Y(n_31) );
AOI221xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_24), .B1(n_27), .B2(n_14), .C(n_28), .Y(n_32) );
AO21x1_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_25), .B(n_5), .Y(n_33) );
AOI221xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_14), .B1(n_25), .B2(n_8), .C(n_1), .Y(n_34) );
UNKNOWN g35 ( );
NAND4xp25_ASAP7_75t_L g36 ( .A(n_32), .B(n_7), .C(n_8), .D(n_14), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
XOR2xp5_ASAP7_75t_L g38 ( .A(n_36), .B(n_14), .Y(n_38) );
BUFx2_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
OAI22x1_ASAP7_75t_SL g40 ( .A1(n_38), .A2(n_35), .B1(n_14), .B2(n_10), .Y(n_40) );
OA22x2_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .B1(n_14), .B2(n_9), .Y(n_41) );
endmodule