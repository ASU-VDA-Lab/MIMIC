module fake_netlist_6_3712_n_1924 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1924);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1924;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVxp33_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_72),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_65),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_110),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_92),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_50),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_24),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_145),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_0),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_32),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_54),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_66),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_54),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_22),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_150),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_120),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_59),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_4),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_22),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_106),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_100),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_2),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_111),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_41),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_93),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_52),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_85),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_155),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_170),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_25),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_177),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_158),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_27),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_127),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_131),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_40),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_98),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_107),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_12),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_52),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_53),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_147),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_68),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_132),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_165),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_80),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_108),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_105),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_172),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_168),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_71),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_28),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_43),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_11),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_97),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_30),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_90),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_6),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_78),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_69),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_64),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_104),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_38),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_182),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_73),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_152),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_124),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_160),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_171),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_34),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_42),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_64),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_68),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_89),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_35),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_154),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_119),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_63),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_70),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_1),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_163),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_77),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_82),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_81),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_137),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_129),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_146),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_75),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_95),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_26),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_62),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_113),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_130),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_142),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_41),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_40),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_180),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_139),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_109),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_88),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_30),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_31),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_118),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_32),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_16),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_15),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_87),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_167),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_91),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_20),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_49),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_13),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_161),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_9),
.Y(n_354)
);

BUFx4f_ASAP7_75t_SL g355 ( 
.A(n_141),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_83),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_148),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_126),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_79),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_39),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_33),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_10),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_66),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_58),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_24),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_112),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_214),
.B(n_3),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_214),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_195),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_203),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_271),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_227),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_229),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_214),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_242),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_214),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_214),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_250),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_239),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_292),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_3),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_202),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_257),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_202),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_185),
.B(n_5),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_240),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_244),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_214),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_214),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_214),
.B(n_5),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_282),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_212),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_276),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_282),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_247),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_282),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_248),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_282),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_282),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_282),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_251),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_191),
.B(n_8),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_200),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_252),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_191),
.B(n_8),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_323),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_282),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_256),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_282),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_255),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_260),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_265),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_236),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_200),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_288),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_197),
.B(n_10),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_211),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_255),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_201),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_211),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_190),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_255),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_204),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_291),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_212),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_255),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_193),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_197),
.B(n_12),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_238),
.B(n_13),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_297),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_189),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_255),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_303),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_293),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_355),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_305),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_207),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_238),
.B(n_14),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_293),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_293),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_293),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_342),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_293),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_204),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_267),
.B(n_317),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_308),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_308),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_308),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_308),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_308),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_208),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_353),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_205),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_264),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_384),
.B(n_186),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_450),
.A2(n_317),
.B(n_267),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_386),
.B(n_186),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_425),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_447),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_394),
.B(n_187),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_387),
.B(n_274),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_425),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_414),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_302),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_425),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_302),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_405),
.B(n_187),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_189),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_376),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_376),
.Y(n_483)
);

AND3x2_ASAP7_75t_L g484 ( 
.A(n_420),
.B(n_328),
.C(n_319),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_423),
.B(n_319),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_378),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_253),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_411),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_427),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_408),
.B(n_325),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_378),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_188),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_437),
.B(n_439),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_439),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_375),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_188),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_390),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_192),
.Y(n_510)
);

XNOR2x2_ASAP7_75t_R g511 ( 
.A(n_371),
.B(n_14),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_391),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_449),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_459),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_382),
.B(n_328),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_391),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_448),
.B(n_253),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_369),
.B(n_321),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_450),
.A2(n_233),
.B(n_208),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_396),
.B(n_211),
.Y(n_523)
);

CKINVDCx6p67_ASAP7_75t_R g524 ( 
.A(n_374),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_380),
.A2(n_254),
.B1(n_198),
.B2(n_262),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_452),
.B(n_453),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_454),
.B(n_192),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_396),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_455),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_418),
.B(n_273),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_383),
.B(n_264),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_369),
.B(n_233),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_474),
.B(n_373),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_463),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_483),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_483),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_469),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_471),
.B(n_381),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_538),
.A2(n_460),
.B1(n_286),
.B2(n_344),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_434),
.C(n_433),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_383),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_476),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_426),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_538),
.A2(n_443),
.B1(n_392),
.B2(n_380),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_492),
.B(n_388),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_492),
.B(n_389),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_462),
.B(n_374),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_515),
.B(n_460),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_489),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_538),
.A2(n_392),
.B1(n_237),
.B2(n_362),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_474),
.B(n_398),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_493),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_502),
.B(n_400),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_469),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_476),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_474),
.B(n_211),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_538),
.A2(n_237),
.B1(n_362),
.B2(n_277),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_538),
.A2(n_277),
.B1(n_334),
.B2(n_273),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_533),
.A2(n_315),
.B1(n_347),
.B2(n_228),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_476),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_502),
.B(n_404),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_534),
.B(n_417),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_499),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_480),
.Y(n_588)
);

INVx4_ASAP7_75t_SL g589 ( 
.A(n_523),
.Y(n_589)
);

BUFx6f_ASAP7_75t_SL g590 ( 
.A(n_502),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_502),
.B(n_407),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_502),
.B(n_412),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_499),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_533),
.B(n_415),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_489),
.B(n_457),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_477),
.B(n_416),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_520),
.B(n_426),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_509),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_419),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_524),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_520),
.A2(n_334),
.B1(n_428),
.B2(n_287),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_478),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_429),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_509),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_519),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_519),
.B(n_456),
.Y(n_609)
);

INVx6_ASAP7_75t_L g610 ( 
.A(n_535),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_432),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_462),
.B(n_435),
.Y(n_612)
);

NOR2x1p5_ASAP7_75t_L g613 ( 
.A(n_524),
.B(n_205),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_536),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_486),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_512),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_465),
.B(n_438),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_512),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_535),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_465),
.B(n_441),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_520),
.A2(n_272),
.B1(n_281),
.B2(n_283),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_516),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_470),
.B(n_451),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_522),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_470),
.B(n_458),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_520),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_463),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_521),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_522),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_467),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_480),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_535),
.B(n_401),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_467),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_535),
.B(n_401),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_478),
.B(n_457),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_520),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_536),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_520),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_482),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_482),
.B(n_402),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_523),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_494),
.B(n_397),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_523),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_473),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_479),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_490),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_479),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_463),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_508),
.A2(n_440),
.B1(n_372),
.B2(n_377),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_484),
.B(n_402),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_463),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_490),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_491),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_482),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_482),
.Y(n_663)
);

NOR3xp33_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_442),
.C(n_432),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_484),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_534),
.B(n_508),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_480),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_514),
.B(n_264),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_480),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_486),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_488),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_514),
.B(n_278),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_482),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_498),
.B(n_211),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_397),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_498),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_481),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_498),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_491),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_503),
.B(n_278),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_498),
.B(n_403),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_498),
.B(n_403),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_505),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_495),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_410),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_505),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_554),
.B(n_488),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_606),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_612),
.B(n_505),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_666),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_556),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_622),
.B(n_505),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_636),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_636),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_626),
.B(n_503),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_629),
.B(n_510),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_657),
.B(n_513),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_558),
.B(n_513),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_576),
.B(n_642),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_556),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_560),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_550),
.B(n_529),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_529),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_550),
.B(n_196),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_575),
.B(n_196),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_675),
.B(n_650),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_568),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_650),
.B(n_481),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_581),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_564),
.B(n_194),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_643),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_605),
.B(n_539),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_605),
.B(n_206),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_609),
.B(n_481),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_643),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_639),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_539),
.B(n_206),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_569),
.B(n_385),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_559),
.B(n_658),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_559),
.B(n_215),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_658),
.B(n_215),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_658),
.B(n_564),
.Y(n_726)
);

NOR2x1p5_ASAP7_75t_L g727 ( 
.A(n_548),
.B(n_524),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_609),
.B(n_572),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_670),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_641),
.B(n_521),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_591),
.A2(n_521),
.B(n_442),
.C(n_341),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_649),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_610),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_609),
.B(n_481),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_563),
.B(n_595),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_572),
.B(n_481),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_641),
.B(n_521),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_553),
.B(n_525),
.C(n_234),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_601),
.B(n_518),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_610),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_610),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_601),
.B(n_518),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_618),
.B(n_615),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_602),
.B(n_395),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_608),
.B(n_216),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_649),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_608),
.B(n_518),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_652),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_652),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_671),
.B(n_496),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_687),
.B(n_518),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_596),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_547),
.B(n_490),
.C(n_241),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_518),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_665),
.B(n_216),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_653),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_646),
.B(n_518),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_665),
.B(n_223),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_642),
.A2(n_409),
.B1(n_356),
.B2(n_357),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_567),
.A2(n_464),
.B1(n_485),
.B2(n_531),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_653),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_655),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_661),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_552),
.A2(n_298),
.B1(n_285),
.B2(n_199),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_518),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_661),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_671),
.B(n_223),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_679),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_685),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_687),
.B(n_662),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_577),
.A2(n_464),
.B1(n_485),
.B2(n_531),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_680),
.B(n_224),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_668),
.B(n_224),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_672),
.B(n_225),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_663),
.B(n_530),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_685),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_663),
.B(n_530),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_673),
.B(n_530),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_573),
.B(n_532),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_676),
.B(n_530),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_552),
.A2(n_225),
.B1(n_226),
.B2(n_310),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_599),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_584),
.B(n_226),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_676),
.B(n_530),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_678),
.B(n_683),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_549),
.A2(n_632),
.B1(n_552),
.B2(n_623),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_678),
.B(n_530),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_590),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_555),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_549),
.A2(n_338),
.B1(n_217),
.B2(n_218),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_596),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_614),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_627),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_552),
.B(n_464),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_683),
.B(n_531),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_542),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_599),
.B(n_485),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_645),
.A2(n_485),
.B1(n_531),
.B2(n_523),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_570),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_542),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_604),
.B(n_592),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_645),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_632),
.A2(n_531),
.B(n_485),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_570),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_593),
.B(n_310),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_571),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_627),
.B(n_531),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_549),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_549),
.A2(n_531),
.B1(n_523),
.B2(n_266),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_632),
.A2(n_497),
.B(n_495),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_638),
.A2(n_640),
.B(n_647),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_543),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_599),
.B(n_497),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_543),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_561),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_585),
.B(n_312),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_630),
.B(n_312),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_561),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_599),
.A2(n_320),
.B1(n_294),
.B2(n_263),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_630),
.B(n_313),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_580),
.A2(n_511),
.B1(n_307),
.B2(n_222),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_571),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_562),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_587),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_681),
.A2(n_501),
.B(n_500),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_610),
.B(n_500),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_587),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_562),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_600),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_630),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_620),
.B(n_501),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_611),
.B(n_313),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_620),
.B(n_504),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_611),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_620),
.B(n_504),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_620),
.B(n_506),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_576),
.B(n_506),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_607),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_576),
.B(n_507),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_576),
.A2(n_523),
.B1(n_210),
.B2(n_231),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_566),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_576),
.B(n_507),
.Y(n_846)
);

INVxp33_ASAP7_75t_L g847 ( 
.A(n_580),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_682),
.B(n_517),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_644),
.B(n_318),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_654),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_611),
.B(n_318),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_689),
.B(n_696),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_733),
.A2(n_686),
.B(n_635),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_806),
.A2(n_617),
.B(n_607),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_691),
.B(n_644),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_697),
.B(n_611),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_704),
.B(n_619),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_688),
.B(n_660),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_708),
.B(n_710),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_544),
.Y(n_861)
);

CKINVDCx10_ASAP7_75t_R g862 ( 
.A(n_824),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_837),
.B(n_613),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_735),
.A2(n_590),
.B1(n_644),
.B2(n_613),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_850),
.B(n_544),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_740),
.A2(n_637),
.B(n_588),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_730),
.A2(n_624),
.B(n_621),
.Y(n_867)
);

AND2x2_ASAP7_75t_SL g868 ( 
.A(n_786),
.B(n_578),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_702),
.B(n_621),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_743),
.B(n_574),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_843),
.B(n_574),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_740),
.A2(n_637),
.B(n_579),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_721),
.B(n_738),
.C(n_744),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_740),
.A2(n_637),
.B(n_579),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_736),
.A2(n_582),
.B(n_566),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_739),
.A2(n_586),
.B(n_582),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_741),
.A2(n_565),
.B(n_555),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_741),
.A2(n_565),
.B(n_555),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_723),
.A2(n_590),
.B1(n_669),
.B2(n_633),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_741),
.A2(n_565),
.B(n_555),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_706),
.B(n_624),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_715),
.A2(n_625),
.B(n_633),
.C(n_594),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_810),
.A2(n_565),
.B(n_555),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_784),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_729),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_706),
.B(n_625),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_742),
.A2(n_594),
.B(n_586),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_747),
.A2(n_616),
.B(n_598),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_709),
.B(n_598),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_784),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_847),
.A2(n_358),
.B(n_349),
.C(n_346),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_760),
.A2(n_628),
.B(n_616),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_709),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_805),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_717),
.A2(n_634),
.B(n_541),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_712),
.B(n_540),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_734),
.A2(n_541),
.B(n_540),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_752),
.B(n_603),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_805),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_781),
.B(n_684),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_714),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_714),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_718),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_718),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_692),
.B(n_540),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_690),
.A2(n_333),
.B1(n_230),
.B2(n_243),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_785),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_711),
.B(n_541),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_693),
.B(n_545),
.Y(n_909)
);

O2A1O1Ixp5_ASAP7_75t_L g910 ( 
.A1(n_703),
.A2(n_804),
.B(n_813),
.C(n_814),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_750),
.B(n_728),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_794),
.B(n_551),
.Y(n_912)
);

OAI22x1_ASAP7_75t_L g913 ( 
.A1(n_727),
.A2(n_307),
.B1(n_306),
.B2(n_314),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_694),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_773),
.A2(n_583),
.B(n_545),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_795),
.B(n_583),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_737),
.B(n_583),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_843),
.B(n_603),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_737),
.A2(n_656),
.B(n_631),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_713),
.B(n_631),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_808),
.B(n_791),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_700),
.A2(n_656),
.B(n_631),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_713),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_726),
.A2(n_527),
.B(n_528),
.C(n_537),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_816),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_694),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_713),
.B(n_656),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_775),
.B(n_259),
.C(n_246),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_700),
.A2(n_659),
.B(n_565),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_719),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_796),
.B(n_589),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_720),
.B(n_232),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_755),
.B(n_331),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_805),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_805),
.B(n_684),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_719),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_695),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_789),
.A2(n_669),
.B1(n_332),
.B2(n_339),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_722),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_722),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_776),
.B(n_232),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_724),
.B(n_232),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_816),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_748),
.B(n_659),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_769),
.B(n_245),
.Y(n_946)
);

AOI33xp33_ASAP7_75t_L g947 ( 
.A1(n_765),
.A2(n_258),
.A3(n_284),
.B1(n_290),
.B2(n_295),
.B3(n_300),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_772),
.A2(n_788),
.B(n_754),
.C(n_757),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_837),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_829),
.A2(n_667),
.B(n_677),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_731),
.A2(n_343),
.B(n_304),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_749),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_749),
.B(n_667),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_833),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_834),
.A2(n_838),
.B(n_836),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_791),
.B(n_331),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_761),
.B(n_667),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_839),
.A2(n_801),
.B(n_766),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_677),
.B(n_684),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_732),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_758),
.B(n_332),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_762),
.B(n_677),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_800),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_732),
.Y(n_964)
);

BUFx4f_ASAP7_75t_L g965 ( 
.A(n_800),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_764),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_745),
.A2(n_725),
.B(n_705),
.C(n_716),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_698),
.B(n_245),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_811),
.A2(n_669),
.B1(n_337),
.B2(n_336),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_SL g970 ( 
.A1(n_777),
.A2(n_363),
.B(n_330),
.C(n_345),
.Y(n_970)
);

NOR2x1_ASAP7_75t_L g971 ( 
.A(n_833),
.B(n_528),
.Y(n_971)
);

NOR2x1_ASAP7_75t_L g972 ( 
.A(n_820),
.B(n_823),
.Y(n_972)
);

NOR2x1p5_ASAP7_75t_SL g973 ( 
.A(n_799),
.B(n_410),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_746),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_759),
.B(n_336),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_811),
.B(n_684),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_797),
.A2(n_767),
.B1(n_768),
.B2(n_778),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_779),
.A2(n_684),
.B(n_557),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_768),
.B(n_537),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_707),
.A2(n_316),
.B(n_322),
.C(n_311),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_780),
.A2(n_684),
.B(n_651),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_783),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_771),
.B(n_337),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_774),
.B(n_245),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_819),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_L g986 ( 
.A1(n_835),
.A2(n_220),
.B(n_213),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_778),
.B(n_339),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_851),
.A2(n_219),
.B(n_209),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_746),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_756),
.A2(n_413),
.B(n_309),
.C(n_361),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_756),
.B(n_360),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_763),
.B(n_360),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_763),
.B(n_361),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_849),
.B(n_368),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_770),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_793),
.B(n_551),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_782),
.A2(n_651),
.B(n_648),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_770),
.B(n_368),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_822),
.A2(n_413),
.B(n_468),
.C(n_461),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_797),
.A2(n_249),
.B1(n_327),
.B2(n_359),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_797),
.A2(n_249),
.B1(n_327),
.B2(n_359),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_802),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_753),
.B(n_209),
.Y(n_1003)
);

AO22x1_ASAP7_75t_L g1004 ( 
.A1(n_792),
.A2(n_306),
.B1(n_219),
.B2(n_220),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_802),
.B(n_674),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_807),
.B(n_674),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_812),
.B(n_551),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_807),
.B(n_674),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_797),
.B(n_840),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_809),
.B(n_825),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_787),
.A2(n_790),
.B(n_798),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_809),
.B(n_589),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_825),
.B(n_674),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_827),
.B(n_589),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_848),
.A2(n_557),
.B(n_651),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_827),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_830),
.B(n_674),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_830),
.B(n_674),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_832),
.B(n_674),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_841),
.A2(n_523),
.B1(n_249),
.B2(n_359),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_842),
.A2(n_651),
.B(n_648),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_832),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_846),
.A2(n_651),
.B(n_648),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_828),
.A2(n_648),
.B(n_557),
.Y(n_1024)
);

OAI321xp33_ASAP7_75t_L g1025 ( 
.A1(n_859),
.A2(n_852),
.A3(n_984),
.B1(n_942),
.B2(n_986),
.C(n_988),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_860),
.B(n_799),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_899),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1002),
.Y(n_1028)
);

AND2x4_ASAP7_75t_SL g1029 ( 
.A(n_954),
.B(n_803),
.Y(n_1029)
);

BUFx4_ASAP7_75t_SL g1030 ( 
.A(n_863),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_885),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_SL g1032 ( 
.A1(n_891),
.A2(n_845),
.B(n_815),
.C(n_831),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1016),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_861),
.B(n_340),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_899),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_856),
.A2(n_845),
.B(n_817),
.C(n_831),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_907),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_871),
.B(n_817),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_857),
.B(n_818),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_868),
.B(n_818),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_866),
.A2(n_844),
.B(n_826),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_940),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_925),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_944),
.B(n_870),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1022),
.B(n_821),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_982),
.B(n_865),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_963),
.B(n_965),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_911),
.B(n_826),
.Y(n_1048)
);

O2A1O1Ixp5_ASAP7_75t_L g1049 ( 
.A1(n_910),
.A2(n_468),
.B(n_461),
.C(n_472),
.Y(n_1049)
);

CKINVDCx14_ASAP7_75t_R g1050 ( 
.A(n_918),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_949),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_967),
.A2(n_472),
.B(n_278),
.C(n_301),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_858),
.A2(n_340),
.B1(n_327),
.B2(n_359),
.Y(n_1053)
);

O2A1O1Ixp5_ASAP7_75t_L g1054 ( 
.A1(n_1000),
.A2(n_472),
.B(n_301),
.C(n_324),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_968),
.B(n_340),
.Y(n_1055)
);

OAI22x1_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_367),
.B1(n_366),
.B2(n_365),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_932),
.B(n_261),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_893),
.B(n_268),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_940),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_975),
.A2(n_994),
.B(n_933),
.C(n_961),
.Y(n_1060)
);

AO22x1_ASAP7_75t_L g1061 ( 
.A1(n_972),
.A2(n_367),
.B1(n_366),
.B2(n_365),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_1010),
.A2(n_327),
.B1(n_359),
.B2(n_324),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_901),
.B(n_269),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_1001),
.A2(n_472),
.B(n_324),
.C(n_301),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_1012),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_902),
.B(n_270),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_977),
.A2(n_327),
.B1(n_279),
.B2(n_280),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1003),
.B(n_275),
.Y(n_1068)
);

AND2x2_ASAP7_75t_SL g1069 ( 
.A(n_963),
.B(n_84),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_289),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_903),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_867),
.A2(n_955),
.B(n_853),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_R g1073 ( 
.A(n_965),
.B(n_213),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_1012),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_884),
.B(n_589),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_985),
.A2(n_296),
.B(n_299),
.C(n_350),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_904),
.B(n_351),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_930),
.B(n_352),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_943),
.B(n_354),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_884),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_936),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_952),
.B(n_326),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_898),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_966),
.B(n_326),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_899),
.A2(n_364),
.B1(n_329),
.B2(n_314),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_934),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_898),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1014),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_863),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_928),
.A2(n_364),
.B(n_329),
.C(n_222),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_906),
.A2(n_221),
.B(n_17),
.C(n_19),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_884),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_946),
.B(n_921),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_990),
.A2(n_221),
.B(n_17),
.C(n_19),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_890),
.B(n_475),
.Y(n_1095)
);

AND2x2_ASAP7_75t_SL g1096 ( 
.A(n_934),
.B(n_184),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_934),
.A2(n_475),
.B1(n_466),
.B2(n_181),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_958),
.A2(n_475),
.B(n_466),
.C(n_21),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_890),
.B(n_15),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_890),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_894),
.B(n_179),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_863),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_917),
.A2(n_475),
.B(n_466),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

OR2x2_ASAP7_75t_SL g1105 ( 
.A(n_862),
.B(n_20),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_960),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_855),
.A2(n_466),
.B1(n_169),
.B2(n_166),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_854),
.A2(n_157),
.B(n_156),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_R g1109 ( 
.A(n_954),
.B(n_136),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_983),
.B(n_21),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_869),
.B(n_23),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_954),
.B(n_134),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_939),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_987),
.B(n_991),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_939),
.B(n_125),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1014),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_958),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_947),
.B(n_29),
.C(n_36),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_894),
.A2(n_121),
.B1(n_116),
.B2(n_103),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_960),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_951),
.A2(n_926),
.B1(n_941),
.B2(n_974),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_971),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_914),
.A2(n_995),
.B1(n_989),
.B2(n_937),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_913),
.A2(n_36),
.B(n_37),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_881),
.B(n_37),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_956),
.B(n_38),
.C(n_43),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1009),
.B(n_931),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_973),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_964),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_886),
.B(n_964),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_889),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_931),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_872),
.A2(n_101),
.B(n_99),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_872),
.A2(n_49),
.B(n_53),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_SL g1135 ( 
.A1(n_938),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_908),
.B(n_1011),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1004),
.B(n_56),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_992),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_SL g1139 ( 
.A(n_969),
.B(n_57),
.C(n_60),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1011),
.B(n_60),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_R g1141 ( 
.A(n_1009),
.B(n_61),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_993),
.B(n_61),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_998),
.B(n_62),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_874),
.A2(n_63),
.B(n_65),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_979),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_1009),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_920),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_927),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_915),
.A2(n_71),
.B1(n_896),
.B2(n_905),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_882),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_980),
.B(n_879),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_909),
.B(n_919),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_919),
.B(n_916),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_915),
.A2(n_897),
.B(n_895),
.C(n_892),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_945),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_924),
.B(n_1020),
.C(n_999),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_953),
.B(n_962),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_957),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_912),
.B(n_948),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_935),
.Y(n_1160)
);

OAI22x1_ASAP7_75t_L g1161 ( 
.A1(n_976),
.A2(n_900),
.B1(n_996),
.B2(n_1007),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1005),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_874),
.A2(n_978),
.B(n_997),
.Y(n_1163)
);

CKINVDCx8_ASAP7_75t_R g1164 ( 
.A(n_970),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1006),
.B(n_1008),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1044),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1034),
.B(n_895),
.Y(n_1167)
);

AO32x2_ASAP7_75t_L g1168 ( 
.A1(n_1149),
.A2(n_875),
.A3(n_876),
.B1(n_888),
.B2(n_887),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1028),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1145),
.B(n_875),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_1013),
.B1(n_1017),
.B2(n_1018),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1060),
.A2(n_1019),
.B1(n_897),
.B2(n_929),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1033),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_1031),
.B(n_929),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1136),
.A2(n_950),
.B(n_883),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1163),
.A2(n_922),
.B(n_878),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1152),
.A2(n_1026),
.B(n_1153),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1025),
.A2(n_887),
.B(n_888),
.C(n_1015),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_1154),
.A2(n_877),
.B(n_880),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1114),
.B(n_959),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_1068),
.A2(n_1015),
.B1(n_959),
.B2(n_1024),
.C(n_1021),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1114),
.B(n_981),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1039),
.A2(n_1023),
.B(n_1157),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1157),
.A2(n_1041),
.B(n_1130),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1048),
.A2(n_1159),
.B(n_1140),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1057),
.B(n_1055),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1131),
.B(n_1040),
.Y(n_1187)
);

CKINVDCx11_ASAP7_75t_R g1188 ( 
.A(n_1037),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1089),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1027),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_R g1191 ( 
.A(n_1050),
.B(n_1080),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1071),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1051),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1081),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1030),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_1103),
.B(n_1108),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1079),
.A2(n_1093),
.B1(n_1138),
.B2(n_1110),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1038),
.B(n_1079),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1165),
.A2(n_1032),
.B(n_1036),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1110),
.A2(n_1052),
.B(n_1151),
.C(n_1142),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1098),
.A2(n_1165),
.B(n_1049),
.Y(n_1201)
);

AOI21xp33_ASAP7_75t_L g1202 ( 
.A1(n_1143),
.A2(n_1111),
.B(n_1125),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1117),
.A2(n_1115),
.B(n_1112),
.C(n_1128),
.Y(n_1203)
);

INVx5_ASAP7_75t_L g1204 ( 
.A(n_1027),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1133),
.A2(n_1047),
.B(n_1155),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_SL g1206 ( 
.A1(n_1076),
.A2(n_1075),
.B(n_1090),
.C(n_1147),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1096),
.B(n_1069),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1121),
.A2(n_1144),
.B(n_1134),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1031),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1082),
.B(n_1084),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1043),
.B(n_1083),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1162),
.A2(n_1097),
.A3(n_1148),
.B(n_1056),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_1067),
.A2(n_1135),
.A3(n_1119),
.B1(n_1085),
.B2(n_1139),
.Y(n_1214)
);

OAI222xp33_ASAP7_75t_L g1215 ( 
.A1(n_1091),
.A2(n_1137),
.B1(n_1062),
.B2(n_1053),
.C1(n_1094),
.C2(n_1043),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_1092),
.B(n_1078),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1054),
.A2(n_1064),
.B(n_1123),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1054),
.A2(n_1064),
.B(n_1156),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1087),
.A2(n_1069),
.B1(n_1122),
.B2(n_1070),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1123),
.A2(n_1129),
.B(n_1062),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1045),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1118),
.A2(n_1107),
.B(n_1066),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1058),
.A2(n_1077),
.B(n_1063),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1096),
.A2(n_1095),
.B(n_1127),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1100),
.B(n_1127),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_SL g1226 ( 
.A1(n_1120),
.A2(n_1059),
.B(n_1106),
.C(n_1042),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1139),
.A2(n_1053),
.B(n_1120),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1099),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1070),
.B(n_1061),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1127),
.A2(n_1146),
.B(n_1029),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1027),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_1116),
.B(n_1074),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1073),
.B(n_1124),
.C(n_1164),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1065),
.B(n_1074),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1141),
.A2(n_1102),
.B1(n_1126),
.B2(n_1146),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1088),
.B(n_1132),
.Y(n_1236)
);

AOI221x1_ASAP7_75t_L g1237 ( 
.A1(n_1099),
.A2(n_1160),
.B1(n_1141),
.B2(n_1113),
.C(n_1086),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1088),
.B(n_1132),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1146),
.A2(n_1160),
.B1(n_1035),
.B2(n_1086),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1146),
.A2(n_1104),
.B(n_1035),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1073),
.Y(n_1241)
);

AO21x1_ASAP7_75t_L g1242 ( 
.A1(n_1101),
.A2(n_1160),
.B(n_1035),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1105),
.A2(n_1030),
.B(n_1109),
.C(n_1101),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1035),
.Y(n_1244)
);

NAND3x1_ASAP7_75t_L g1245 ( 
.A(n_1086),
.B(n_1104),
.C(n_1113),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1104),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1113),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1154),
.A2(n_1072),
.A3(n_1098),
.B(n_1159),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1051),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_SL g1250 ( 
.A1(n_1140),
.A2(n_689),
.B(n_1001),
.C(n_1000),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1034),
.B(n_870),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1060),
.B(n_852),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1154),
.A2(n_1072),
.A3(n_1098),
.B(n_1159),
.Y(n_1253)
);

OAI21xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1062),
.A2(n_689),
.B(n_852),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1060),
.A2(n_689),
.B(n_1117),
.C(n_804),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1031),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1037),
.Y(n_1257)
);

INVx6_ASAP7_75t_L g1258 ( 
.A(n_1037),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1132),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1072),
.A2(n_740),
.B(n_733),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1060),
.B(n_852),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1037),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1060),
.A2(n_689),
.B1(n_852),
.B2(n_1062),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1060),
.B(n_852),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1080),
.B(n_1100),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1072),
.A2(n_740),
.B(n_733),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1027),
.Y(n_1267)
);

AOI22x1_ASAP7_75t_L g1268 ( 
.A1(n_1161),
.A2(n_1150),
.B1(n_1151),
.B2(n_984),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1154),
.A2(n_1072),
.A3(n_1098),
.B(n_1159),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1060),
.A2(n_689),
.B(n_910),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_SL g1271 ( 
.A1(n_1060),
.A2(n_689),
.B(n_1117),
.C(n_804),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_SL g1272 ( 
.A(n_1060),
.B(n_689),
.C(n_873),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_1099),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1154),
.A2(n_1072),
.A3(n_1098),
.B(n_1159),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1060),
.A2(n_689),
.B(n_859),
.C(n_852),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1034),
.B(n_870),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1060),
.A2(n_689),
.B(n_852),
.C(n_873),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1028),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1037),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1060),
.A2(n_689),
.B(n_852),
.C(n_873),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1046),
.B(n_689),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1037),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1051),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1060),
.A2(n_689),
.B(n_859),
.C(n_852),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1060),
.A2(n_689),
.B(n_910),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1037),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1034),
.B(n_870),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1060),
.B(n_852),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1145),
.B(n_852),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1072),
.A2(n_1154),
.B(n_1163),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1060),
.A2(n_847),
.B1(n_859),
.B2(n_699),
.C(n_688),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1072),
.A2(n_1154),
.B(n_1163),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1060),
.A2(n_689),
.B(n_852),
.C(n_873),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_R g1294 ( 
.A(n_1050),
.B(n_544),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1028),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1051),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1072),
.A2(n_1154),
.B(n_1163),
.Y(n_1297)
);

INVx3_ASAP7_75t_SL g1298 ( 
.A(n_1089),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1060),
.A2(n_847),
.B1(n_859),
.B2(n_699),
.C(n_688),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1060),
.A2(n_689),
.B(n_852),
.C(n_873),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1068),
.A2(n_689),
.B1(n_868),
.B2(n_847),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1145),
.B(n_852),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1028),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1060),
.A2(n_740),
.B(n_733),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1145),
.B(n_852),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1145),
.B(n_852),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1060),
.B(n_870),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1060),
.A2(n_689),
.B(n_852),
.C(n_873),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1145),
.B(n_852),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1173),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_1301),
.B2(n_1198),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1241),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1272),
.A2(n_1307),
.B1(n_1261),
.B2(n_1288),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1252),
.A2(n_1264),
.B1(n_1263),
.B2(n_1229),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1188),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1192),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1258),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1207),
.A2(n_1263),
.B1(n_1281),
.B2(n_1251),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1289),
.B(n_1302),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1207),
.A2(n_1276),
.B1(n_1287),
.B2(n_1273),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1309),
.B1(n_1306),
.B2(n_1305),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1294),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1258),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1295),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1211),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1233),
.A2(n_1222),
.B1(n_1202),
.B2(n_1254),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1289),
.A2(n_1309),
.B1(n_1306),
.B2(n_1305),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1262),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1204),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1279),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1222),
.A2(n_1202),
.B1(n_1285),
.B2(n_1270),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1169),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1177),
.A2(n_1266),
.B(n_1260),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1302),
.A2(n_1219),
.B1(n_1228),
.B2(n_1200),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1204),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1270),
.A2(n_1285),
.B1(n_1210),
.B2(n_1223),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1194),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1223),
.A2(n_1227),
.B1(n_1268),
.B2(n_1167),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1236),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1227),
.A2(n_1218),
.B1(n_1235),
.B2(n_1273),
.Y(n_1341)
);

INVx8_ASAP7_75t_L g1342 ( 
.A(n_1204),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1191),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1187),
.B(n_1221),
.Y(n_1344)
);

BUFx4f_ASAP7_75t_SL g1345 ( 
.A(n_1189),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1218),
.A2(n_1180),
.B1(n_1166),
.B2(n_1187),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1278),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1303),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1180),
.A2(n_1166),
.B1(n_1182),
.B2(n_1186),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1259),
.Y(n_1350)
);

INVx6_ASAP7_75t_L g1351 ( 
.A(n_1267),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1275),
.B(n_1284),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1211),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1225),
.B(n_1265),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1236),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1231),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1257),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1216),
.A2(n_1308),
.B1(n_1300),
.B2(n_1277),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1298),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1248),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1237),
.A2(n_1212),
.B1(n_1256),
.B2(n_1170),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1174),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1282),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1267),
.B(n_1239),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1170),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1280),
.B(n_1293),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1286),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1209),
.Y(n_1368)
);

BUFx4f_ASAP7_75t_SL g1369 ( 
.A(n_1265),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1224),
.A2(n_1236),
.B1(n_1234),
.B2(n_1172),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1234),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1226),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1193),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1249),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1232),
.Y(n_1375)
);

BUFx4_ASAP7_75t_R g1376 ( 
.A(n_1243),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1248),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1297),
.A2(n_1201),
.B1(n_1208),
.B2(n_1290),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1171),
.A2(n_1242),
.B1(n_1225),
.B2(n_1181),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1267),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1246),
.Y(n_1381)
);

BUFx2_ASAP7_75t_SL g1382 ( 
.A(n_1190),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1238),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1283),
.B(n_1296),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1190),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1247),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1201),
.A2(n_1208),
.B1(n_1292),
.B2(n_1290),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1255),
.A2(n_1271),
.B1(n_1206),
.B2(n_1203),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1292),
.A2(n_1185),
.B1(n_1184),
.B2(n_1217),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1217),
.A2(n_1215),
.B1(n_1220),
.B2(n_1230),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1183),
.A2(n_1205),
.B1(n_1220),
.B2(n_1199),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1304),
.A2(n_1178),
.B1(n_1245),
.B2(n_1240),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1179),
.A2(n_1214),
.B1(n_1176),
.B2(n_1175),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1244),
.A2(n_1214),
.B1(n_1213),
.B2(n_1250),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_SL g1395 ( 
.A(n_1213),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1213),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1214),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1248),
.A2(n_1274),
.B1(n_1269),
.B2(n_1253),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1168),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1253),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1196),
.A2(n_1269),
.B1(n_1274),
.B2(n_1168),
.Y(n_1403)
);

BUFx8_ASAP7_75t_L g1404 ( 
.A(n_1168),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1274),
.A2(n_1299),
.B1(n_1291),
.B2(n_689),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1207),
.A2(n_689),
.B1(n_1198),
.B2(n_847),
.Y(n_1406)
);

CKINVDCx6p67_ASAP7_75t_R g1407 ( 
.A(n_1188),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1258),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1207),
.A2(n_689),
.B1(n_1229),
.B2(n_859),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1258),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1411)
);

INVx8_ASAP7_75t_L g1412 ( 
.A(n_1204),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1173),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1188),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1258),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1173),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1188),
.Y(n_1417)
);

CKINVDCx6p67_ASAP7_75t_R g1418 ( 
.A(n_1188),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1204),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1173),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1258),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1204),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1207),
.A2(n_689),
.B1(n_1198),
.B2(n_847),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1188),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1427)
);

CKINVDCx16_ASAP7_75t_R g1428 ( 
.A(n_1294),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1291),
.A2(n_689),
.B1(n_1060),
.B2(n_859),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1173),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1173),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1291),
.A2(n_689),
.B1(n_1060),
.B2(n_859),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1207),
.A2(n_689),
.B1(n_1229),
.B2(n_859),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1251),
.B(n_1276),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1258),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1188),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1204),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1207),
.A2(n_689),
.B1(n_1198),
.B2(n_847),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1188),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1262),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1198),
.B(n_852),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1258),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1211),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1173),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_689),
.B2(n_1301),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1258),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1258),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1399),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1402),
.B(n_1325),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1335),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1319),
.B(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1360),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1333),
.A2(n_1389),
.B(n_1391),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1311),
.A2(n_1429),
.B1(n_1432),
.B2(n_1411),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1404),
.A2(n_1400),
.B1(n_1334),
.B2(n_1397),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1377),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1321),
.B(n_1344),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1371),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1401),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1404),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1389),
.A2(n_1391),
.B(n_1403),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1398),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1364),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1353),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1442),
.B(n_1325),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1398),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1411),
.A2(n_1427),
.B1(n_1423),
.B2(n_1424),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1375),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1395),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1395),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1444),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1365),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1335),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1353),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1368),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1409),
.B(n_1433),
.Y(n_1479)
);

AO31x2_ASAP7_75t_L g1480 ( 
.A1(n_1394),
.A2(n_1352),
.A3(n_1392),
.B(n_1366),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1364),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1396),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1332),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1338),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1372),
.A2(n_1362),
.B(n_1348),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1393),
.A2(n_1387),
.B(n_1378),
.Y(n_1486)
);

AND2x2_ASAP7_75t_SL g1487 ( 
.A(n_1378),
.B(n_1387),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1347),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1310),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1370),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1335),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1316),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1370),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1349),
.B(n_1423),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1417),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1324),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1358),
.B(n_1350),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1388),
.A2(n_1331),
.B(n_1313),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1413),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1416),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1331),
.A2(n_1313),
.B(n_1339),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1420),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1342),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1430),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1336),
.B(n_1314),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1431),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1445),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1336),
.B(n_1314),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1381),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1339),
.A2(n_1326),
.B(n_1379),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1426),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1346),
.B(n_1326),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1434),
.Y(n_1515)
);

BUFx8_ASAP7_75t_L g1516 ( 
.A(n_1414),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1356),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_SL g1518 ( 
.A(n_1312),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1351),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1390),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1383),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1342),
.B(n_1412),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1405),
.A2(n_1341),
.B(n_1346),
.Y(n_1523)
);

AOI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1424),
.A2(n_1446),
.B(n_1441),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1342),
.B(n_1412),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1361),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1361),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1349),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1427),
.A2(n_1446),
.B1(n_1441),
.B2(n_1318),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1436),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1406),
.A2(n_1425),
.B(n_1438),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1341),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1405),
.B(n_1406),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1412),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1384),
.A2(n_1437),
.B(n_1351),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1351),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1437),
.A2(n_1380),
.B(n_1419),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1425),
.Y(n_1539)
);

NAND2x1_ASAP7_75t_L g1540 ( 
.A(n_1380),
.B(n_1419),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1438),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1320),
.B(n_1354),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1329),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1329),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1374),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1422),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1354),
.A2(n_1357),
.B1(n_1428),
.B2(n_1386),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1376),
.A2(n_1382),
.B(n_1385),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1312),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1369),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1328),
.B(n_1440),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1369),
.A2(n_1373),
.B(n_1363),
.Y(n_1552)
);

AOI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1323),
.A2(n_1415),
.B(n_1317),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1448),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1448),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1317),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1330),
.B(n_1367),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1317),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1455),
.A2(n_1524),
.B(n_1470),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1477),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1552),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1462),
.B(n_1410),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1462),
.B(n_1408),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1542),
.B(n_1408),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_R g1565 ( 
.A(n_1530),
.B(n_1315),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1452),
.B(n_1447),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1529),
.A2(n_1418),
.B1(n_1407),
.B2(n_1343),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1479),
.A2(n_1359),
.B1(n_1322),
.B2(n_1345),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1485),
.A2(n_1345),
.B(n_1421),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1466),
.B(n_1439),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1477),
.B(n_1421),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_SL g1573 ( 
.A(n_1474),
.B(n_1337),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1483),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_L g1575 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_SL g1576 ( 
.A1(n_1482),
.A2(n_1435),
.B(n_1443),
.C(n_1447),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1512),
.A2(n_1435),
.B(n_1443),
.C(n_1447),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1474),
.B(n_1435),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1532),
.A2(n_1527),
.B(n_1533),
.C(n_1495),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1467),
.B(n_1490),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1503),
.A2(n_1500),
.B(n_1523),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1553),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1523),
.A2(n_1500),
.B(n_1491),
.C(n_1494),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_SL g1584 ( 
.A(n_1522),
.B(n_1525),
.Y(n_1584)
);

OAI211xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1547),
.A2(n_1526),
.B(n_1555),
.C(n_1554),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1491),
.A2(n_1494),
.B(n_1527),
.C(n_1514),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_SL g1587 ( 
.A1(n_1482),
.A2(n_1468),
.B(n_1532),
.C(n_1478),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1507),
.A2(n_1510),
.B(n_1533),
.Y(n_1588)
);

NAND2x1_ASAP7_75t_L g1589 ( 
.A(n_1522),
.B(n_1525),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1507),
.A2(n_1510),
.B(n_1514),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1558),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1521),
.Y(n_1592)
);

AO32x2_ASAP7_75t_L g1593 ( 
.A1(n_1451),
.A2(n_1519),
.A3(n_1537),
.B1(n_1476),
.B2(n_1492),
.Y(n_1593)
);

AO32x1_ASAP7_75t_L g1594 ( 
.A1(n_1526),
.A2(n_1520),
.A3(n_1461),
.B1(n_1459),
.B2(n_1453),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_R g1595 ( 
.A(n_1550),
.B(n_1557),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1456),
.A2(n_1520),
.B(n_1541),
.C(n_1539),
.Y(n_1596)
);

AO32x2_ASAP7_75t_L g1597 ( 
.A1(n_1451),
.A2(n_1519),
.A3(n_1492),
.B1(n_1476),
.B2(n_1537),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1539),
.A2(n_1541),
.B(n_1528),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1547),
.A2(n_1481),
.B(n_1465),
.C(n_1528),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1499),
.A2(n_1531),
.B1(n_1550),
.B2(n_1465),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1496),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1511),
.B(n_1499),
.C(n_1545),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1558),
.A2(n_1531),
.B(n_1555),
.C(n_1554),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1558),
.Y(n_1604)
);

AND2x4_ASAP7_75t_SL g1605 ( 
.A(n_1557),
.B(n_1496),
.Y(n_1605)
);

INVx4_ASAP7_75t_SL g1606 ( 
.A(n_1536),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_SL g1607 ( 
.A(n_1549),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1465),
.B(n_1481),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1499),
.A2(n_1486),
.B(n_1487),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1513),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1481),
.B(n_1472),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1475),
.B(n_1460),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_SL g1613 ( 
.A1(n_1540),
.A2(n_1473),
.B(n_1472),
.C(n_1550),
.Y(n_1613)
);

AND2x2_ASAP7_75t_SL g1614 ( 
.A(n_1499),
.B(n_1487),
.Y(n_1614)
);

OAI211xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1501),
.A2(n_1509),
.B(n_1508),
.C(n_1506),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1487),
.A2(n_1548),
.B(n_1535),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1548),
.A2(n_1553),
.B(n_1538),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1549),
.Y(n_1618)
);

AO21x2_ASAP7_75t_L g1619 ( 
.A1(n_1449),
.A2(n_1464),
.B(n_1469),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1489),
.B(n_1493),
.Y(n_1620)
);

BUFx12f_ASAP7_75t_L g1621 ( 
.A(n_1513),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1469),
.A2(n_1531),
.B1(n_1498),
.B2(n_1502),
.C(n_1504),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1484),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1473),
.B(n_1489),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1460),
.B(n_1480),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1493),
.B(n_1497),
.Y(n_1626)
);

NAND4xp25_ASAP7_75t_L g1627 ( 
.A(n_1549),
.B(n_1509),
.C(n_1502),
.D(n_1504),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1609),
.B(n_1454),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1574),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1626),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1609),
.B(n_1454),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1626),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1559),
.A2(n_1463),
.B1(n_1516),
.B2(n_1498),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1623),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1586),
.A2(n_1450),
.B1(n_1488),
.B2(n_1463),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1620),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1463),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1457),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1559),
.A2(n_1450),
.B1(n_1488),
.B2(n_1518),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1625),
.B(n_1457),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1612),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1619),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1560),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1621),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1606),
.Y(n_1646)
);

AND4x1_ASAP7_75t_L g1647 ( 
.A(n_1579),
.B(n_1543),
.C(n_1546),
.D(n_1544),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1449),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1589),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1584),
.B(n_1471),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1593),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1594),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1594),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1594),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1597),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1480),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1602),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1608),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1634),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1634),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1651),
.B(n_1602),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1633),
.A2(n_1614),
.B1(n_1575),
.B2(n_1588),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1643),
.A2(n_1617),
.B(n_1570),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1660),
.A2(n_1590),
.B1(n_1588),
.B2(n_1603),
.C(n_1583),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1643),
.A2(n_1617),
.B(n_1577),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1650),
.B(n_1608),
.Y(n_1669)
);

INVx5_ASAP7_75t_SL g1670 ( 
.A(n_1652),
.Y(n_1670)
);

OAI322xp33_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1567),
.A3(n_1578),
.B1(n_1572),
.B2(n_1600),
.C1(n_1568),
.C2(n_1604),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1580),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1633),
.A2(n_1596),
.B1(n_1590),
.B2(n_1585),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1640),
.A2(n_1595),
.B1(n_1567),
.B2(n_1599),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1660),
.A2(n_1587),
.B1(n_1598),
.B2(n_1576),
.C(n_1627),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1644),
.Y(n_1676)
);

BUFx2_ASAP7_75t_SL g1677 ( 
.A(n_1646),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1635),
.A2(n_1613),
.B(n_1582),
.C(n_1550),
.Y(n_1678)
);

OAI33xp33_ASAP7_75t_L g1679 ( 
.A1(n_1651),
.A2(n_1627),
.A3(n_1506),
.B1(n_1501),
.B2(n_1508),
.B3(n_1517),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1660),
.A2(n_1569),
.B1(n_1571),
.B2(n_1598),
.C(n_1618),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1635),
.A2(n_1573),
.B1(n_1564),
.B2(n_1607),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1638),
.B(n_1592),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1644),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1661),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1630),
.B(n_1566),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1636),
.B(n_1624),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1639),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1639),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1640),
.A2(n_1591),
.B(n_1611),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1629),
.Y(n_1693)
);

NAND4xp25_ASAP7_75t_L g1694 ( 
.A(n_1651),
.B(n_1561),
.C(n_1563),
.D(n_1562),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1629),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1652),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1629),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1639),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1641),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1641),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1693),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1686),
.B(n_1689),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1693),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1695),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_R g1709 ( 
.A(n_1687),
.B(n_1601),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1698),
.B(n_1696),
.Y(n_1711)
);

NAND2x1p5_ASAP7_75t_L g1712 ( 
.A(n_1664),
.B(n_1647),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1686),
.B(n_1649),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1695),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1667),
.A2(n_1628),
.B1(n_1631),
.B2(n_1635),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1698),
.B(n_1649),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1696),
.B(n_1649),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1697),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1663),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1686),
.B(n_1653),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1670),
.B(n_1661),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1683),
.B(n_1642),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1701),
.B(n_1653),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_L g1729 ( 
.A(n_1664),
.B(n_1646),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1662),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1701),
.B(n_1654),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1689),
.B(n_1654),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1701),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1662),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1702),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1701),
.B(n_1654),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1670),
.B(n_1658),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1663),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1663),
.Y(n_1741)
);

OAI32xp33_ASAP7_75t_L g1742 ( 
.A1(n_1680),
.A2(n_1659),
.A3(n_1658),
.B1(n_1640),
.B2(n_1657),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1742),
.B(n_1645),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1712),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1712),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1704),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1728),
.B(n_1689),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1706),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1715),
.A2(n_1681),
.B1(n_1673),
.B2(n_1665),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1670),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1742),
.B(n_1645),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1712),
.B(n_1690),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1669),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1735),
.B(n_1685),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1669),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1737),
.B(n_1669),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1717),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1708),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1708),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1729),
.B(n_1685),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1714),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1729),
.B(n_1675),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1707),
.B(n_1690),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1707),
.B(n_1690),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1737),
.B(n_1646),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1717),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1714),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1722),
.B(n_1648),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1738),
.A2(n_1673),
.B1(n_1674),
.B2(n_1665),
.Y(n_1772)
);

NAND2x1_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1658),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1718),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1678),
.C(n_1674),
.D(n_1692),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1722),
.B(n_1699),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1725),
.B(n_1648),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1717),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1718),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1727),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1669),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1647),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1727),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1725),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1730),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1756),
.B(n_1758),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1758),
.B(n_1711),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1765),
.B(n_1699),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_SL g1791 ( 
.A(n_1775),
.B(n_1645),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1757),
.B(n_1682),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.B(n_1677),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1751),
.B(n_1699),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1772),
.B(n_1688),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1753),
.B(n_1700),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1773),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1763),
.B(n_1688),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1744),
.B(n_1645),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1773),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1745),
.B(n_1700),
.Y(n_1801)
);

AO22x1_ASAP7_75t_L g1802 ( 
.A1(n_1785),
.A2(n_1516),
.B1(n_1610),
.B2(n_1740),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1782),
.B(n_1677),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1770),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1782),
.B(n_1700),
.Y(n_1805)
);

NAND2x1_ASAP7_75t_L g1806 ( 
.A(n_1752),
.B(n_1733),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1746),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1752),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1755),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1746),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1705),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1747),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1755),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1747),
.Y(n_1814)
);

NAND2x1_ASAP7_75t_L g1815 ( 
.A(n_1759),
.B(n_1733),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1782),
.B(n_1647),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1749),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1756),
.B(n_1648),
.Y(n_1818)
);

NAND2x1_ASAP7_75t_L g1819 ( 
.A(n_1759),
.B(n_1733),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1750),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1761),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1754),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1781),
.B(n_1703),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1784),
.B(n_1648),
.Y(n_1824)
);

OAI332xp33_ASAP7_75t_L g1825 ( 
.A1(n_1816),
.A2(n_1754),
.A3(n_1769),
.B1(n_1760),
.B2(n_1778),
.B3(n_1768),
.C1(n_1659),
.C2(n_1777),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1807),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1802),
.A2(n_1671),
.B(n_1668),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1791),
.A2(n_1709),
.B(n_1781),
.C(n_1628),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1793),
.A2(n_1668),
.B(n_1762),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1799),
.A2(n_1637),
.B1(n_1631),
.B2(n_1628),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1810),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1794),
.B(n_1795),
.Y(n_1833)
);

O2A1O1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1804),
.A2(n_1764),
.B(n_1783),
.C(n_1780),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1808),
.B(n_1787),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1812),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1808),
.A2(n_1787),
.B1(n_1631),
.B2(n_1628),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1814),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1817),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1799),
.B(n_1516),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_L g1841 ( 
.A(n_1822),
.B(n_1679),
.C(n_1774),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1822),
.B(n_1779),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1796),
.A2(n_1668),
.B(n_1786),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1788),
.A2(n_1637),
.B1(n_1631),
.B2(n_1668),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1820),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1803),
.A2(n_1806),
.B(n_1790),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1792),
.B(n_1516),
.Y(n_1847)
);

NOR4xp25_ASAP7_75t_L g1848 ( 
.A(n_1809),
.B(n_1813),
.C(n_1821),
.D(n_1805),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_L g1849 ( 
.A(n_1809),
.B(n_1769),
.C(n_1760),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1813),
.A2(n_1643),
.B1(n_1710),
.B2(n_1703),
.C(n_1716),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1832),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1833),
.A2(n_1803),
.B1(n_1788),
.B2(n_1789),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1828),
.A2(n_1803),
.B1(n_1819),
.B2(n_1815),
.Y(n_1853)
);

OAI32xp33_ASAP7_75t_L g1854 ( 
.A1(n_1841),
.A2(n_1800),
.A3(n_1797),
.B1(n_1824),
.B2(n_1658),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1847),
.B(n_1823),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1848),
.A2(n_1801),
.B(n_1800),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1840),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1826),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1835),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1827),
.A2(n_1789),
.B1(n_1823),
.B2(n_1637),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1831),
.Y(n_1861)
);

AOI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1834),
.A2(n_1798),
.B(n_1797),
.Y(n_1862)
);

NOR3xp33_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1811),
.C(n_1818),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1836),
.Y(n_1864)
);

O2A1O1Ixp33_ASAP7_75t_SL g1865 ( 
.A1(n_1846),
.A2(n_1565),
.B(n_1658),
.C(n_1650),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1838),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1846),
.A2(n_1605),
.B(n_1766),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1843),
.B(n_1666),
.C(n_1766),
.Y(n_1868)
);

OAI211xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1829),
.A2(n_1778),
.B(n_1776),
.C(n_1767),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1839),
.Y(n_1870)
);

O2A1O1Ixp33_ASAP7_75t_SL g1871 ( 
.A1(n_1854),
.A2(n_1842),
.B(n_1845),
.C(n_1850),
.Y(n_1871)
);

OAI32xp33_ASAP7_75t_L g1872 ( 
.A1(n_1863),
.A2(n_1849),
.A3(n_1837),
.B1(n_1850),
.B2(n_1716),
.Y(n_1872)
);

OAI221xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1852),
.A2(n_1844),
.B1(n_1830),
.B2(n_1748),
.C(n_1767),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1851),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1866),
.B(n_1851),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1853),
.A2(n_1650),
.B1(n_1637),
.B2(n_1666),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1866),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1855),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1857),
.A2(n_1552),
.B(n_1776),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1856),
.B(n_1666),
.C(n_1748),
.Y(n_1881)
);

NOR4xp25_ASAP7_75t_L g1882 ( 
.A(n_1871),
.B(n_1870),
.C(n_1858),
.D(n_1861),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1875),
.Y(n_1883)
);

NOR3x1_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1864),
.C(n_1868),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1879),
.B(n_1859),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1878),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1878),
.B(n_1855),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1881),
.B(n_1860),
.C(n_1857),
.Y(n_1888)
);

NOR2xp67_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1867),
.Y(n_1889)
);

NAND2x1_ASAP7_75t_L g1890 ( 
.A(n_1877),
.B(n_1865),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_L g1891 ( 
.A(n_1873),
.B(n_1862),
.C(n_1869),
.Y(n_1891)
);

AOI222xp33_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_1872),
.B1(n_1854),
.B2(n_1865),
.C1(n_1876),
.C2(n_1710),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1882),
.A2(n_1710),
.B1(n_1716),
.B2(n_1726),
.C(n_1711),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1890),
.A2(n_1740),
.B(n_1726),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1887),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_SL g1896 ( 
.A(n_1888),
.B(n_1684),
.C(n_1711),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1883),
.A2(n_1719),
.B1(n_1724),
.B2(n_1736),
.C(n_1731),
.Y(n_1897)
);

NOR4xp25_ASAP7_75t_L g1898 ( 
.A(n_1886),
.B(n_1731),
.C(n_1719),
.D(n_1736),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1895),
.A2(n_1885),
.B(n_1884),
.C(n_1889),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1896),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1894),
.B(n_1893),
.Y(n_1901)
);

OAI322xp33_ASAP7_75t_L g1902 ( 
.A1(n_1892),
.A2(n_1721),
.A3(n_1713),
.B1(n_1732),
.B2(n_1657),
.C1(n_1655),
.C2(n_1656),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1898),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1897),
.A2(n_1726),
.B1(n_1724),
.B2(n_1736),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1903),
.B(n_1900),
.Y(n_1905)
);

NAND2xp33_ASAP7_75t_L g1906 ( 
.A(n_1899),
.B(n_1902),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1901),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1904),
.A2(n_1726),
.B1(n_1719),
.B2(n_1724),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1900),
.Y(n_1909)
);

NOR3xp33_ASAP7_75t_L g1910 ( 
.A(n_1907),
.B(n_1646),
.C(n_1540),
.Y(n_1910)
);

NOR2xp67_ASAP7_75t_L g1911 ( 
.A(n_1909),
.B(n_1713),
.Y(n_1911)
);

NOR3xp33_ASAP7_75t_L g1912 ( 
.A(n_1905),
.B(n_1906),
.C(n_1908),
.Y(n_1912)
);

AND2x2_ASAP7_75t_SL g1913 ( 
.A(n_1912),
.B(n_1646),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1913),
.A2(n_1910),
.B1(n_1911),
.B2(n_1726),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1914),
.B(n_1731),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1914),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1916),
.B(n_1721),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1915),
.Y(n_1918)
);

OA21x2_ASAP7_75t_L g1919 ( 
.A1(n_1917),
.A2(n_1720),
.B(n_1741),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1919),
.B(n_1918),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1732),
.B(n_1705),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1921),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_R g1923 ( 
.A1(n_1922),
.A2(n_1741),
.B1(n_1720),
.B2(n_1666),
.C(n_1734),
.Y(n_1923)
);

AOI211xp5_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1534),
.B(n_1505),
.C(n_1536),
.Y(n_1924)
);


endmodule