module fake_jpeg_15512_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_8),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_20),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_56),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_71),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_81),
.B1(n_24),
.B2(n_31),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_63),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_29),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_29),
.B1(n_28),
.B2(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_29),
.B1(n_28),
.B2(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_28),
.B1(n_16),
.B2(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_62),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_20),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_102)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_22),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_51),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_31),
.B(n_22),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_48),
.B(n_56),
.C(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_24),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_121),
.B1(n_125),
.B2(n_78),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_55),
.A3(n_39),
.B1(n_37),
.B2(n_61),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_71),
.A3(n_79),
.B1(n_76),
.B2(n_46),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_61),
.B1(n_52),
.B2(n_57),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_117),
.B1(n_69),
.B2(n_78),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_66),
.C(n_60),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_110),
.C(n_115),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_21),
.B(n_23),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_33),
.B(n_18),
.C(n_32),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_118),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_66),
.C(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_52),
.B1(n_58),
.B2(n_51),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_0),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_1),
.B(n_2),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_52),
.B1(n_58),
.B2(n_51),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_86),
.C(n_76),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_122),
.C(n_123),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_137),
.B1(n_141),
.B2(n_150),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_80),
.B1(n_82),
.B2(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_140),
.B1(n_146),
.B2(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_89),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_104),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_149),
.B(n_27),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_142),
.B(n_143),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_97),
.B1(n_70),
.B2(n_69),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_70),
.B1(n_84),
.B2(n_46),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_1),
.B(n_2),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_123),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_99),
.A2(n_76),
.B1(n_71),
.B2(n_32),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

NOR2x1p5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_46),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_66),
.B1(n_91),
.B2(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_137),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_169),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_108),
.A3(n_101),
.B1(n_117),
.B2(n_124),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_172),
.B1(n_174),
.B2(n_112),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_159),
.B(n_162),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_101),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_171),
.C(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_R g161 ( 
.A(n_149),
.B(n_102),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_177),
.B(n_142),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_148),
.B(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_135),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_145),
.B1(n_138),
.B2(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_107),
.B1(n_103),
.B2(n_125),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_129),
.B1(n_127),
.B2(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_105),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_122),
.A3(n_33),
.B1(n_18),
.B2(n_32),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_98),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_135),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_128),
.C(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_183),
.B1(n_195),
.B2(n_204),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_131),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_188),
.C(n_196),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_191),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_134),
.B(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_187),
.B1(n_194),
.B2(n_197),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_144),
.C(n_150),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_141),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_158),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_203),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_163),
.B1(n_161),
.B2(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_130),
.B1(n_140),
.B2(n_134),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_134),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_171),
.B1(n_153),
.B2(n_166),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_112),
.B1(n_91),
.B2(n_98),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_116),
.B1(n_18),
.B2(n_27),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_98),
.B1(n_119),
.B2(n_32),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_155),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_206),
.B(n_217),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_165),
.B1(n_159),
.B2(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_225),
.B1(n_202),
.B2(n_23),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_162),
.C(n_158),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_228),
.C(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_156),
.B1(n_170),
.B2(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_227),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_177),
.C(n_173),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_186),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_184),
.B(n_185),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_236),
.B1(n_241),
.B2(n_247),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_197),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_218),
.C(n_219),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_201),
.B1(n_186),
.B2(n_188),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_216),
.B1(n_237),
.B2(n_249),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_183),
.B1(n_178),
.B2(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_170),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_226),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_192),
.B1(n_179),
.B2(n_172),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_26),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_119),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_2),
.B(n_3),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_23),
.B1(n_21),
.B2(n_5),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_260),
.C(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_26),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_216),
.B1(n_208),
.B2(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_258),
.B1(n_270),
.B2(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_210),
.B1(n_227),
.B2(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_218),
.C(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_265),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_224),
.C(n_213),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_221),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_269),
.C(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_213),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_119),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_17),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_250),
.B(n_247),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_235),
.C(n_236),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_119),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_231),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_275),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_245),
.C(n_251),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_250),
.B1(n_251),
.B2(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_279),
.A2(n_263),
.B1(n_252),
.B2(n_26),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_14),
.B1(n_4),
.B2(n_6),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_26),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_284),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_14),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_3),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_278),
.B1(n_276),
.B2(n_271),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_290),
.B1(n_300),
.B2(n_9),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_258),
.B(n_254),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_273),
.B(n_8),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_255),
.B1(n_257),
.B2(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_7),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_273),
.B1(n_284),
.B2(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_304),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_26),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_17),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_8),
.C(n_9),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_9),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_10),
.B(n_11),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_9),
.B(n_10),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_10),
.Y(n_311)
);

AOI21x1_ASAP7_75t_SL g312 ( 
.A1(n_288),
.A2(n_10),
.B(n_11),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_300),
.C(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_314),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_290),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_297),
.B(n_293),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_297),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_320),
.B(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_327),
.B1(n_11),
.B2(n_12),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_320),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_315),
.B(n_12),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_330),
.B1(n_322),
.B2(n_326),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_12),
.B(n_13),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_13),
.C(n_331),
.Y(n_335)
);


endmodule