module fake_jpeg_16461_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_56),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_34),
.B1(n_19),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_50),
.B1(n_55),
.B2(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_18),
.B2(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_20),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_17),
.B(n_33),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_17),
.B(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_32),
.B1(n_22),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_88),
.B1(n_89),
.B2(n_23),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_35),
.Y(n_113)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_34),
.B(n_15),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_91),
.Y(n_98)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_SL g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_22),
.B1(n_23),
.B2(n_30),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_124),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_0),
.B(n_1),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_45),
.C(n_43),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_121),
.C(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_34),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_54),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_25),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_35),
.B1(n_86),
.B2(n_74),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_120),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_24),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_45),
.C(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_67),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_125),
.B(n_124),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_115),
.B1(n_122),
.B2(n_130),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_70),
.B(n_97),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_155),
.B(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_73),
.B1(n_76),
.B2(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_97),
.B1(n_76),
.B2(n_70),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_143),
.B1(n_153),
.B2(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_103),
.B1(n_110),
.B2(n_77),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_80),
.B1(n_75),
.B2(n_93),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_29),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_150),
.B(n_110),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_105),
.C(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_98),
.A2(n_80),
.B1(n_75),
.B2(n_52),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_111),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_95),
.B1(n_77),
.B2(n_26),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_176),
.C(n_146),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_182),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_165),
.B1(n_155),
.B2(n_154),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_170),
.B(n_171),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_123),
.B1(n_119),
.B2(n_106),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_174),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_119),
.B1(n_106),
.B2(n_120),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_99),
.B1(n_104),
.B2(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_95),
.B1(n_102),
.B2(n_14),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_115),
.B1(n_102),
.B2(n_26),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_128),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_102),
.B1(n_13),
.B2(n_15),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_185),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_115),
.B1(n_117),
.B2(n_25),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_184),
.B(n_24),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_29),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

XOR2x2_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_24),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_137),
.B1(n_129),
.B2(n_140),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_24),
.B1(n_21),
.B2(n_2),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_168),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_192),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_127),
.B1(n_141),
.B2(n_153),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_196),
.B1(n_205),
.B2(n_216),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_139),
.B(n_138),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_197),
.B(n_200),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_198),
.C(n_206),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_143),
.B1(n_152),
.B2(n_130),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_145),
.C(n_25),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_145),
.B1(n_28),
.B2(n_21),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_10),
.B(n_15),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_14),
.C(n_13),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_94),
.Y(n_202)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_172),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_117),
.B(n_28),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_21),
.C(n_24),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_158),
.B1(n_175),
.B2(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_0),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_1),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_161),
.B1(n_184),
.B2(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_220),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_242),
.B1(n_199),
.B2(n_197),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_208),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_167),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_229),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_196),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_160),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_182),
.C(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_237),
.C(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_190),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_234),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_239),
.B1(n_227),
.B2(n_205),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_189),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_194),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_172),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_180),
.B1(n_174),
.B2(n_177),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_245),
.A2(n_235),
.B1(n_221),
.B2(n_200),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_251),
.B1(n_266),
.B2(n_205),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_242),
.B1(n_227),
.B2(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_204),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_260),
.B(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_206),
.C(n_210),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_225),
.C(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_193),
.B(n_178),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_210),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_212),
.B1(n_193),
.B2(n_205),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_240),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_229),
.C(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_221),
.C(n_191),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_279),
.B1(n_249),
.B2(n_247),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_244),
.B(n_254),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_193),
.B1(n_226),
.B2(n_213),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_170),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_181),
.C(n_3),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_2),
.Y(n_298)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_260),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_285),
.B(n_273),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_258),
.C(n_253),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_249),
.B(n_252),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_292),
.B1(n_295),
.B2(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_256),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_283),
.B(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_296),
.C(n_270),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_263),
.B1(n_282),
.B2(n_284),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_3),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_301),
.C(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_267),
.C(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_261),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_308),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_4),
.C(n_5),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_5),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_289),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_288),
.C(n_295),
.Y(n_315)
);

AOI21x1_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_310),
.B(n_300),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_285),
.B(n_290),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_290),
.B(n_12),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_10),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_301),
.C(n_305),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_323),
.A2(n_329),
.B(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_325),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_314),
.C(n_322),
.Y(n_330)
);

AO21x1_ASAP7_75t_SL g329 ( 
.A1(n_313),
.A2(n_11),
.B(n_7),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_332),
.A3(n_328),
.B1(n_326),
.B2(n_333),
.C(n_9),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_6),
.B(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_7),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_8),
.B1(n_9),
.B2(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);


endmodule