module fake_jpeg_23838_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_22),
.B(n_30),
.C(n_25),
.Y(n_56)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_49),
.B1(n_41),
.B2(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_19),
.B1(n_32),
.B2(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_22),
.B(n_25),
.C(n_24),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_92)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_75),
.B(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_78),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_89),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_35),
.B(n_17),
.C(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_87),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_39),
.C(n_40),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_91),
.C(n_22),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_57),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_27),
.B1(n_17),
.B2(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_33),
.Y(n_98)
);

OR2x4_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_22),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_22),
.B(n_40),
.C(n_36),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_102),
.B(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_90),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_47),
.B1(n_63),
.B2(n_52),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_47),
.B1(n_40),
.B2(n_61),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_109),
.B1(n_115),
.B2(n_117),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_47),
.B1(n_40),
.B2(n_17),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_96),
.B1(n_70),
.B2(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_80),
.B1(n_67),
.B2(n_70),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_85),
.C(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_24),
.B1(n_23),
.B2(n_21),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_39),
.B(n_22),
.C(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_100),
.C(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_130),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_116),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_145),
.B(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_73),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_71),
.B1(n_95),
.B2(n_103),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_153),
.B1(n_103),
.B2(n_21),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_144),
.B(n_90),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_83),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_79),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_79),
.A3(n_93),
.B1(n_66),
.B2(n_78),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_74),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_119),
.C(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_102),
.B1(n_106),
.B2(n_70),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_168),
.B1(n_133),
.B2(n_152),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_119),
.B(n_120),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_159),
.B(n_170),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_121),
.B1(n_100),
.B2(n_111),
.C(n_125),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_169),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_10),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_121),
.C(n_95),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_93),
.B(n_21),
.C(n_105),
.D(n_125),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_130),
.B(n_128),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

NAND4xp25_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_145),
.C(n_151),
.D(n_143),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_74),
.C(n_16),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_2),
.C(n_3),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_177),
.B(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_127),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_193),
.B1(n_195),
.B2(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_141),
.Y(n_190)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_132),
.B1(n_153),
.B2(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_196),
.B1(n_156),
.B2(n_160),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_142),
.B1(n_149),
.B2(n_150),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_12),
.C(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_135),
.B1(n_145),
.B2(n_131),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_170),
.A3(n_175),
.B1(n_166),
.B2(n_160),
.C1(n_178),
.C2(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_161),
.C(n_165),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_202),
.C(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_171),
.C(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_212),
.B1(n_192),
.B2(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_6),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_208),
.Y(n_225)
);

OAI322xp33_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_191),
.B1(n_194),
.B2(n_181),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_14),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_14),
.C(n_15),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_180),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_196),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_201),
.B(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

AOI31xp67_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_195),
.A3(n_186),
.B(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_220),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_190),
.B1(n_183),
.B2(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_212),
.B1(n_207),
.B2(n_214),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_193),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_223),
.B(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_200),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_233),
.C(n_180),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_215),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_202),
.C(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_210),
.B1(n_193),
.B2(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_240),
.B(n_243),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_225),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_233),
.B(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_247),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_236),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

AOI221xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_251),
.B1(n_232),
.B2(n_221),
.C(n_193),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_252),
.A2(n_228),
.B(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_250),
.Y(n_256)
);


endmodule