module fake_jpeg_5516_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_37),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_44),
.B(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_40),
.B1(n_17),
.B2(n_21),
.Y(n_70)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_20),
.A2(n_10),
.B(n_15),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_56),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_19),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_9),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_36),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_23),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_14),
.Y(n_98)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_71),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_73),
.B(n_81),
.Y(n_129)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_84),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_47),
.B1(n_59),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_77),
.A2(n_80),
.B1(n_91),
.B2(n_32),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_56),
.B1(n_29),
.B2(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_89),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_21),
.B1(n_34),
.B2(n_37),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_14),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_14),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_87),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_24),
.B1(n_36),
.B2(n_33),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_121),
.B1(n_142),
.B2(n_11),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_30),
.B1(n_33),
.B2(n_24),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_119),
.Y(n_162)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_139),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_30),
.B1(n_27),
.B2(n_31),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_30),
.B1(n_31),
.B2(n_6),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_143),
.B(n_32),
.Y(n_165)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_127),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_31),
.B1(n_63),
.B2(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_140),
.B1(n_141),
.B2(n_145),
.Y(n_160)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_113),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_1),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_75),
.B1(n_79),
.B2(n_104),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_73),
.A2(n_64),
.B1(n_63),
.B2(n_60),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_102),
.B1(n_89),
.B2(n_104),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_32),
.Y(n_161)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_76),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_150),
.B(n_170),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_70),
.B(n_81),
.C(n_88),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_79),
.B1(n_83),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_156),
.B1(n_126),
.B2(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_152),
.B(n_164),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_100),
.B(n_97),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_127),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_157),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_64),
.B1(n_108),
.B2(n_109),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_11),
.C(n_16),
.Y(n_157)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_177),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_108),
.B1(n_32),
.B2(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_172),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_1),
.C(n_2),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_175),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_2),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_3),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_128),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_164),
.B1(n_149),
.B2(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_3),
.C(n_5),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_117),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_113),
.B(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_180),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_124),
.B1(n_126),
.B2(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_13),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_214),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_201),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_165),
.B(n_156),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_161),
.B1(n_150),
.B2(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_141),
.B1(n_123),
.B2(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_123),
.B1(n_116),
.B2(n_119),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_133),
.B(n_116),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_163),
.B1(n_166),
.B2(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_203),
.Y(n_221)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_210),
.B1(n_182),
.B2(n_199),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_151),
.A2(n_125),
.B1(n_134),
.B2(n_135),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_212),
.B1(n_175),
.B2(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_167),
.Y(n_218)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_13),
.B1(n_179),
.B2(n_148),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_153),
.C(n_156),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_228),
.C(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_222),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_207),
.B(n_187),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_234),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_155),
.B(n_168),
.C(n_170),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_183),
.B1(n_195),
.B2(n_187),
.Y(n_246)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_173),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_189),
.B(n_183),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_184),
.B1(n_214),
.B2(n_208),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_158),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_158),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_239),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_246),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_257),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_224),
.B(n_216),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_189),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_259),
.C(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_255),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_247),
.B(n_249),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_185),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_202),
.A3(n_197),
.B1(n_188),
.B2(n_201),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_213),
.B(n_203),
.C(n_190),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_218),
.B(n_221),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_190),
.C(n_191),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_268),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_266),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_276),
.B(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_228),
.C(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_215),
.C(n_220),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_242),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_216),
.B1(n_226),
.B2(n_219),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_280)
);

XNOR2x2_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_224),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_287),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_282),
.B(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_268),
.C(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_288),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_258),
.B(n_240),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_246),
.B1(n_261),
.B2(n_271),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_252),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_295),
.B(n_296),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_250),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_269),
.C(n_263),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_261),
.B1(n_271),
.B2(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_299),
.B1(n_285),
.B2(n_280),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_263),
.B1(n_257),
.B2(n_253),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_281),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_302),
.B(n_303),
.Y(n_309)
);

NAND4xp25_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_225),
.C(n_288),
.D(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_248),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_280),
.B(n_224),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_307),
.B(n_250),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_274),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_313),
.Y(n_315)
);

AOI31xp67_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_292),
.A3(n_233),
.B(n_296),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_295),
.Y(n_314)
);

OAI321xp33_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_217),
.A3(n_232),
.B1(n_222),
.B2(n_241),
.C(n_210),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_291),
.C(n_318),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_315),
.Y(n_321)
);


endmodule