module fake_jpeg_4853_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_47),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_20),
.B1(n_17),
.B2(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_33),
.C(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_58),
.B(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_41),
.B1(n_36),
.B2(n_20),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_72),
.B1(n_75),
.B2(n_25),
.Y(n_96)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_41),
.B1(n_17),
.B2(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_26),
.B1(n_31),
.B2(n_16),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_73),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_23),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_24),
.B1(n_36),
.B2(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_18),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_16),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_34),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_94),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_15),
.B(n_31),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_88),
.C(n_102),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_18),
.C(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_81),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_35),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_75),
.B1(n_64),
.B2(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_25),
.B1(n_27),
.B2(n_19),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_16),
.C(n_25),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_73),
.C(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_39),
.B1(n_37),
.B2(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_114),
.B1(n_92),
.B2(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_117),
.B1(n_121),
.B2(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_74),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_35),
.C(n_19),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_27),
.B1(n_35),
.B2(n_19),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_61),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_86),
.B(n_88),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_90),
.A3(n_101),
.B1(n_102),
.B2(n_94),
.C1(n_84),
.C2(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_92),
.B1(n_97),
.B2(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_137),
.B1(n_119),
.B2(n_110),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_98),
.B(n_57),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_120),
.B(n_111),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_115),
.C(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_19),
.B1(n_7),
.B2(n_8),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_136),
.C(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_144),
.B(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_0),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_4),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_2),
.C(n_3),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_149),
.C(n_137),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_7),
.C(n_13),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_2),
.C(n_3),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_133),
.C(n_135),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_128),
.B(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_148),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_154),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_151),
.B(n_5),
.C(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_130),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_161),
.B(n_164),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_141),
.B1(n_144),
.B2(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_153),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_148),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_14),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_12),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_150),
.C(n_146),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_161),
.B(n_10),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_173),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_4),
.B(n_6),
.C(n_10),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_167),
.CI(n_174),
.CON(n_177),
.SN(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_177),
.Y(n_179)
);


endmodule