module fake_jpeg_30180_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx11_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_10),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_51),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_R g85 ( 
.A(n_78),
.B(n_57),
.Y(n_85)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_20),
.C(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_70),
.B1(n_58),
.B2(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_70),
.B1(n_50),
.B2(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_92),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_R g103 ( 
.A(n_85),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_66),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_50),
.B1(n_79),
.B2(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_57),
.B1(n_69),
.B2(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_57),
.Y(n_100)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_61),
.B1(n_68),
.B2(n_71),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_64),
.B(n_62),
.C(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_102),
.B1(n_107),
.B2(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_113),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_59),
.B1(n_23),
.B2(n_24),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_7),
.C(n_8),
.Y(n_129)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_109),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_5),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_9),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_123),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_94),
.B(n_81),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_129),
.B(n_130),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_81),
.B(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_8),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_139),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_124),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_129),
.A3(n_125),
.B1(n_41),
.B2(n_42),
.C1(n_38),
.C2(n_34),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_16),
.B1(n_17),
.B2(n_31),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_147),
.B(n_130),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_48),
.B(n_36),
.C(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_153),
.C(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_116),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_138),
.C(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_119),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_152),
.B(n_155),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_143),
.B(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_149),
.B(n_147),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_131),
.A3(n_134),
.B1(n_142),
.B2(n_145),
.C1(n_147),
.C2(n_155),
.Y(n_162)
);


endmodule