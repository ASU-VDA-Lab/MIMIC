module fake_jpeg_10998_n_650 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_21),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_28),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_60),
.B(n_71),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_65),
.Y(n_131)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_62),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_1),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_76),
.B(n_83),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_1),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_89),
.Y(n_180)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_95),
.Y(n_215)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_107),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_100),
.B(n_52),
.Y(n_186)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_2),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_46),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_116),
.Y(n_151)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_26),
.B(n_2),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_46),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_122),
.Y(n_154)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_35),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_35),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_130),
.B(n_145),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_136),
.B(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_137),
.B(n_149),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_42),
.B1(n_54),
.B2(n_57),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_144),
.A2(n_93),
.B1(n_88),
.B2(n_81),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_26),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_34),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_157),
.B(n_170),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_42),
.B1(n_58),
.B2(n_43),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_160),
.A2(n_177),
.B1(n_63),
.B2(n_114),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_70),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_167),
.B(n_186),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_92),
.B(n_47),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_58),
.B1(n_43),
.B2(n_51),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_178),
.B(n_191),
.Y(n_286)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx12_ASAP7_75t_R g298 ( 
.A(n_187),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_47),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_188),
.B(n_190),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_52),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_70),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_34),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_84),
.B(n_36),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_195),
.B(n_196),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_77),
.B(n_36),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_69),
.A2(n_72),
.B1(n_87),
.B2(n_90),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_118),
.B(n_111),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_77),
.B(n_37),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_205),
.B(n_206),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_51),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_85),
.B(n_37),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_208),
.B(n_209),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_129),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_95),
.B(n_57),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_218),
.Y(n_293)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_53),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_11),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_123),
.B(n_53),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_62),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_219),
.B(n_221),
.Y(n_295)
);

HAxp5_ASAP7_75t_SL g220 ( 
.A(n_64),
.B(n_54),
.CON(n_220),
.SN(n_220)
);

OR2x2_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_2),
.Y(n_244)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_263),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_143),
.B(n_98),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_226),
.Y(n_314)
);

INVx5_ASAP7_75t_SL g227 ( 
.A(n_183),
.Y(n_227)
);

INVx4_ASAP7_75t_SL g328 ( 
.A(n_227),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_229),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_139),
.Y(n_230)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_R g232 ( 
.A(n_131),
.B(n_39),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_232),
.B(n_268),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_177),
.A2(n_39),
.B1(n_33),
.B2(n_112),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_234),
.Y(n_359)
);

OA22x2_ASAP7_75t_L g313 ( 
.A1(n_236),
.A2(n_266),
.B1(n_202),
.B2(n_184),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_160),
.A2(n_201),
.B1(n_152),
.B2(n_141),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_237),
.A2(n_278),
.B1(n_200),
.B2(n_184),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_165),
.B(n_98),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_244),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_243),
.Y(n_354)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_91),
.B1(n_104),
.B2(n_102),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_253),
.A2(n_260),
.B1(n_264),
.B2(n_279),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_254),
.A2(n_259),
.B1(n_197),
.B2(n_174),
.Y(n_356)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_255),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_146),
.B(n_127),
.C(n_80),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_256),
.B(n_185),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_199),
.A2(n_68),
.B1(n_176),
.B2(n_150),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_257),
.A2(n_258),
.B1(n_289),
.B2(n_236),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_176),
.A2(n_150),
.B1(n_164),
.B2(n_193),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_144),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_180),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_180),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_154),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_271),
.Y(n_308)
);

AOI22x1_ASAP7_75t_L g266 ( 
.A1(n_164),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_172),
.A2(n_8),
.B(n_10),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_158),
.Y(n_269)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_158),
.Y(n_270)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_275),
.B(n_291),
.Y(n_311)
);

BUFx4f_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_276),
.Y(n_307)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_179),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_280),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_140),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_168),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_198),
.A2(n_15),
.B(n_16),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_299),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_151),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_155),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_288),
.Y(n_349)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_168),
.A2(n_203),
.B1(n_210),
.B2(n_204),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_294),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_16),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_148),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_296),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_148),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_221),
.Y(n_355)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_159),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_315),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_335),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_222),
.B(n_140),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_331),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_344),
.B1(n_346),
.B2(n_256),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_254),
.A2(n_173),
.B1(n_147),
.B2(n_175),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_330),
.A2(n_356),
.B1(n_278),
.B2(n_229),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_226),
.A2(n_163),
.B(n_132),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_291),
.B(n_247),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_292),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_245),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_204),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_340),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_223),
.B(n_173),
.Y(n_340)
);

OA22x2_ASAP7_75t_SL g342 ( 
.A1(n_244),
.A2(n_147),
.B1(n_134),
.B2(n_185),
.Y(n_342)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_275),
.B(n_174),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_343),
.B(n_347),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_243),
.A2(n_202),
.B1(n_217),
.B2(n_171),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_237),
.A2(n_171),
.B1(n_217),
.B2(n_181),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_197),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_239),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_355),
.B(n_271),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_239),
.B(n_134),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_358),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_360),
.B(n_366),
.C(n_384),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_309),
.B(n_251),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_368),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_362),
.A2(n_367),
.B1(n_314),
.B2(n_322),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_364),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_226),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_273),
.B1(n_281),
.B2(n_241),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_308),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_232),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_372),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_317),
.Y(n_372)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_373),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_312),
.A2(n_234),
.B1(n_263),
.B2(n_132),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_379),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_311),
.B(n_235),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_266),
.B(n_255),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_387),
.B(n_358),
.Y(n_421)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_SL g384 ( 
.A(n_302),
.B(n_224),
.C(n_234),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_340),
.B(n_238),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_396),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_249),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_395),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_392),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_393),
.A2(n_312),
.B1(n_354),
.B2(n_358),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_248),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_394),
.Y(n_428)
);

INVx11_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_306),
.B(n_284),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_399),
.Y(n_415)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_301),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_401),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_317),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_403),
.Y(n_436)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_406),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_228),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_407),
.A2(n_430),
.B1(n_431),
.B2(n_433),
.Y(n_479)
);

OAI32xp33_ASAP7_75t_L g408 ( 
.A1(n_398),
.A2(n_343),
.A3(n_315),
.B1(n_347),
.B2(n_314),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_432),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_429),
.B1(n_435),
.B2(n_440),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_362),
.A2(n_356),
.B1(n_313),
.B2(n_342),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_378),
.A2(n_398),
.B1(n_393),
.B2(n_405),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_313),
.B1(n_302),
.B2(n_342),
.Y(n_431)
);

OAI32xp33_ASAP7_75t_L g432 ( 
.A1(n_374),
.A2(n_352),
.A3(n_310),
.B1(n_313),
.B2(n_351),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_302),
.B1(n_321),
.B2(n_329),
.Y(n_433)
);

OAI32xp33_ASAP7_75t_L g434 ( 
.A1(n_374),
.A2(n_405),
.A3(n_381),
.B1(n_386),
.B2(n_361),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_277),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_367),
.A2(n_349),
.B1(n_329),
.B2(n_305),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_365),
.A2(n_321),
.B(n_333),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_381),
.A2(n_305),
.B1(n_357),
.B2(n_181),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_365),
.A2(n_321),
.B1(n_357),
.B2(n_320),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_404),
.B1(n_385),
.B2(n_307),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_425),
.B(n_376),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_447),
.B(n_452),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_360),
.B1(n_387),
.B2(n_366),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_448),
.A2(n_460),
.B1(n_468),
.B2(n_471),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_371),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g487 ( 
.A1(n_449),
.A2(n_457),
.B(n_461),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_382),
.B1(n_402),
.B2(n_372),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_450),
.A2(n_470),
.B1(n_436),
.B2(n_412),
.Y(n_495)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_440),
.Y(n_451)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_451),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_380),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_401),
.C(n_387),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_456),
.C(n_458),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_467),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_363),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_SL g457 ( 
.A(n_410),
.B(n_384),
.C(n_387),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_400),
.C(n_303),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_303),
.C(n_336),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_436),
.C(n_411),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_413),
.A2(n_369),
.B1(n_370),
.B2(n_395),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_425),
.B(n_334),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_475),
.B1(n_417),
.B2(n_442),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_389),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_427),
.Y(n_464)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_383),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_465),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_396),
.Y(n_467)
);

INVx13_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

BUFx5_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_431),
.A2(n_320),
.B1(n_288),
.B2(n_262),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_435),
.A2(n_388),
.B1(n_391),
.B2(n_390),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_316),
.Y(n_472)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_416),
.A2(n_263),
.B1(n_324),
.B2(n_325),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_473),
.A2(n_418),
.B(n_415),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_414),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_478),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_421),
.A2(n_324),
.B(n_373),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_477),
.A2(n_480),
.B(n_481),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_423),
.B(n_345),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_420),
.A2(n_379),
.B(n_325),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_407),
.A2(n_246),
.B(n_399),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_424),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_483),
.B(n_494),
.Y(n_517)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_458),
.B(n_433),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_491),
.B(n_454),
.Y(n_526)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_493),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_438),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_495),
.A2(n_498),
.B1(n_515),
.B2(n_513),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_509),
.C(n_474),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_455),
.B(n_426),
.Y(n_499)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_499),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_428),
.Y(n_500)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_446),
.A2(n_432),
.B1(n_408),
.B2(n_441),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_502),
.A2(n_470),
.B1(n_462),
.B2(n_467),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_466),
.A2(n_415),
.B(n_444),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_503),
.A2(n_511),
.B(n_485),
.Y(n_542)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_444),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_446),
.Y(n_528)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_510),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_474),
.B(n_466),
.C(n_459),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_428),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_511),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_479),
.A2(n_409),
.B1(n_418),
.B2(n_411),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_513),
.A2(n_442),
.B1(n_422),
.B2(n_417),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_468),
.B(n_414),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_443),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_516),
.B(n_532),
.C(n_534),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_454),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_518),
.B(n_522),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_457),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_530),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_508),
.B(n_486),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_526),
.B(n_544),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_528),
.B(n_540),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_529),
.A2(n_536),
.B1(n_527),
.B2(n_497),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_450),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_500),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_531),
.B(n_539),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_477),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_481),
.C(n_460),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_482),
.A2(n_473),
.B1(n_449),
.B2(n_480),
.Y(n_535)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_535),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_422),
.C(n_445),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_543),
.C(n_545),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_496),
.B(n_482),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_505),
.B(n_419),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_499),
.B(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_541),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_542),
.A2(n_501),
.B(n_498),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_509),
.B(n_443),
.C(n_336),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_503),
.B(n_514),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_550),
.A2(n_557),
.B1(n_561),
.B2(n_562),
.Y(n_571)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_541),
.Y(n_551)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_551),
.Y(n_589)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_525),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_558),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_484),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_554),
.B(n_569),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_527),
.A2(n_502),
.B1(n_504),
.B2(n_507),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_519),
.A2(n_512),
.B1(n_489),
.B2(n_488),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_524),
.A2(n_512),
.B1(n_488),
.B2(n_493),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_563),
.A2(n_469),
.B1(n_484),
.B2(n_419),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_534),
.A2(n_485),
.B1(n_495),
.B2(n_487),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_564),
.A2(n_526),
.B1(n_536),
.B2(n_419),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_542),
.A2(n_501),
.B(n_506),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_568),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_510),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_566),
.Y(n_577)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_521),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_570),
.B(n_318),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_516),
.C(n_530),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_573),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_556),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_559),
.A2(n_533),
.B1(n_537),
.B2(n_528),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_574),
.B(n_560),
.Y(n_605)
);

BUFx24_ASAP7_75t_SL g575 ( 
.A(n_546),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_579),
.Y(n_600)
);

BUFx12f_ASAP7_75t_SL g576 ( 
.A(n_567),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_576),
.A2(n_585),
.B(n_580),
.Y(n_598)
);

INVx13_ASAP7_75t_L g578 ( 
.A(n_566),
.Y(n_578)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_555),
.B(n_517),
.C(n_520),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_517),
.C(n_544),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_545),
.C(n_532),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_562),
.Y(n_584)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_584),
.Y(n_596)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_548),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_587),
.B(n_588),
.Y(n_595)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_590),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_586),
.A2(n_565),
.B(n_549),
.Y(n_591)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_591),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_547),
.C(n_564),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_594),
.B(n_601),
.Y(n_619)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_579),
.B(n_547),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_550),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_602),
.B(n_603),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_560),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_574),
.B(n_563),
.C(n_557),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_604),
.B(n_606),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_605),
.A2(n_587),
.B1(n_571),
.B2(n_577),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_571),
.B(n_561),
.C(n_337),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_581),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_576),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_618),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_611),
.B(n_614),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_591),
.A2(n_584),
.B1(n_577),
.B2(n_589),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_612),
.A2(n_318),
.B1(n_299),
.B2(n_261),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_589),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_600),
.B(n_588),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_616),
.B(n_252),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_578),
.B(n_590),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_617),
.A2(n_620),
.B(n_599),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_337),
.C(n_403),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_596),
.A2(n_592),
.B(n_605),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_602),
.B(n_327),
.C(n_345),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_621),
.B(n_296),
.C(n_287),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_623),
.A2(n_626),
.B(n_632),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_609),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_624),
.A2(n_618),
.B1(n_619),
.B2(n_612),
.Y(n_634)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_615),
.A2(n_595),
.B1(n_606),
.B2(n_593),
.C(n_298),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_621),
.B(n_595),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_627),
.B(n_628),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g629 ( 
.A(n_617),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_630),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_631),
.A2(n_269),
.B(n_280),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_610),
.A2(n_240),
.B(n_270),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_634),
.A2(n_638),
.B(n_230),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_624),
.B(n_613),
.C(n_620),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_635),
.A2(n_636),
.B(n_627),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_622),
.A2(n_608),
.B(n_625),
.Y(n_636)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_640),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_633),
.A2(n_630),
.B(n_242),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_641),
.B(n_642),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_637),
.A2(n_231),
.B(n_276),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_644),
.B(n_639),
.Y(n_646)
);

OAI31xp33_ASAP7_75t_SL g647 ( 
.A1(n_646),
.A2(n_643),
.A3(n_276),
.B(n_163),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_163),
.C(n_161),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_169),
.C(n_16),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_169),
.Y(n_650)
);


endmodule