module fake_jpeg_6437_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_41),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_49),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_52),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_55),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_32),
.B(n_30),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_31),
.B1(n_19),
.B2(n_30),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_31),
.B1(n_37),
.B2(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_31),
.B1(n_37),
.B2(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_84),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_34),
.B1(n_22),
.B2(n_37),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_35),
.C(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_39),
.B1(n_40),
.B2(n_16),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_17),
.B1(n_16),
.B2(n_20),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_58),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_61),
.B(n_41),
.C(n_45),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_81),
.B(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_38),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_49),
.B1(n_66),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_84),
.B1(n_85),
.B2(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_35),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_118),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_110),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_17),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_38),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_20),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_39),
.C(n_81),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_104),
.C(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_131),
.B1(n_142),
.B2(n_148),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_38),
.C(n_89),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_111),
.C(n_89),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_1),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_136),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

BUFx16f_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_85),
.B1(n_68),
.B2(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_92),
.C(n_21),
.Y(n_172)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_59),
.B1(n_51),
.B2(n_38),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_99),
.B1(n_106),
.B2(n_96),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_153),
.B1(n_161),
.B2(n_169),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_158),
.C(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_105),
.B1(n_95),
.B2(n_119),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_111),
.C(n_112),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_113),
.B1(n_115),
.B2(n_114),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_70),
.B(n_92),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_171),
.B(n_172),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_122),
.C(n_123),
.D(n_10),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_117),
.B1(n_80),
.B2(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_174),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_92),
.B(n_21),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_80),
.B1(n_27),
.B2(n_23),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_131),
.B1(n_148),
.B2(n_133),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_21),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_171),
.B(n_142),
.CI(n_138),
.CON(n_182),
.SN(n_182)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_183),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_147),
.B1(n_146),
.B2(n_129),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_172),
.B1(n_164),
.B2(n_18),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_147),
.B(n_129),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_192),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_125),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_141),
.B1(n_122),
.B2(n_123),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_151),
.B1(n_170),
.B2(n_165),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_28),
.B(n_21),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_136),
.C(n_143),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_145),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_194),
.B1(n_182),
.B2(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_211),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_169),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_227),
.B(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_160),
.B1(n_152),
.B2(n_166),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_216),
.B1(n_219),
.B2(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_221),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_136),
.B1(n_134),
.B2(n_107),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_70),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_136),
.B1(n_33),
.B2(n_27),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_33),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_183),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_27),
.B(n_26),
.C(n_23),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_190),
.C(n_201),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_235),
.C(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_247),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_213),
.C(n_205),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_192),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_224),
.C(n_214),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_182),
.B1(n_193),
.B2(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_187),
.C(n_180),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_223),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_187),
.B1(n_178),
.B2(n_199),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_26),
.B1(n_28),
.B2(n_8),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_209),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_216),
.C(n_219),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_214),
.C(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_263),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.C(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_225),
.C(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_226),
.C(n_28),
.Y(n_258)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_28),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_26),
.C(n_23),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_265),
.C(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_7),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_249),
.C(n_230),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_246),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_234),
.B1(n_248),
.B2(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_2),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_276),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_279),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_239),
.C(n_238),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_266),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_255),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_8),
.B1(n_13),
.B2(n_4),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_283),
.Y(n_294)
);

AOI31xp33_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_259),
.A3(n_263),
.B(n_251),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_269),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_260),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_277),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_10),
.B(n_13),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_2),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_301),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_278),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_299),
.B(n_5),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_274),
.B(n_269),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_270),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_270),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_294),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_306),
.B1(n_296),
.B2(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_5),
.C(n_6),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_286),
.C(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_303),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_308),
.B(n_314),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.A3(n_315),
.B1(n_317),
.B2(n_318),
.C1(n_15),
.C2(n_12),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_307),
.B(n_11),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_12),
.C(n_15),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_2),
.C(n_3),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_3),
.C(n_319),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_3),
.Y(n_326)
);


endmodule