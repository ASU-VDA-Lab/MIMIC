module real_aes_16589_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_884;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_880;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_637;
wire n_526;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g897 ( .A(n_0), .B(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_1), .A2(n_34), .B1(n_150), .B2(n_200), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_2), .A2(n_95), .B1(n_121), .B2(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_3), .A2(n_119), .B1(n_120), .B2(n_123), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_3), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_4), .A2(n_11), .B1(n_533), .B2(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g898 ( .A(n_5), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_6), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_7), .A2(n_12), .B1(n_553), .B2(n_554), .Y(n_552) );
OR2x2_ASAP7_75t_L g116 ( .A(n_8), .B(n_30), .Y(n_116) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_9), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_10), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_13), .B(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_14), .A2(n_101), .B1(n_244), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_15), .A2(n_31), .B1(n_564), .B2(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_16), .B(n_165), .Y(n_580) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_17), .A2(n_47), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_18), .B(n_259), .Y(n_258) );
AOI21xp33_ASAP7_75t_L g852 ( .A1(n_19), .A2(n_853), .B(n_860), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_20), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_21), .A2(n_38), .B1(n_220), .B2(n_249), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_22), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_23), .A2(n_44), .B1(n_220), .B2(n_533), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_24), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_25), .B(n_564), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_26), .B(n_194), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_27), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_28), .B(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_29), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_32), .A2(n_85), .B1(n_150), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_33), .A2(n_37), .B1(n_150), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_35), .A2(n_51), .B1(n_533), .B2(n_535), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_36), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_39), .Y(n_869) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_40), .B(n_165), .Y(n_233) );
INVx2_ASAP7_75t_L g111 ( .A(n_41), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_42), .B(n_237), .Y(n_254) );
BUFx3_ASAP7_75t_L g114 ( .A(n_43), .Y(n_114) );
INVx1_ASAP7_75t_L g868 ( .A(n_43), .Y(n_868) );
OAI22x1_ASAP7_75t_SL g874 ( .A1(n_45), .A2(n_875), .B1(n_876), .B2(n_879), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_45), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_46), .B(n_183), .Y(n_261) );
AND2x2_ASAP7_75t_L g222 ( .A(n_48), .B(n_183), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_49), .B(n_180), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_50), .A2(n_81), .B1(n_877), .B2(n_878), .Y(n_876) );
INVxp67_ASAP7_75t_L g877 ( .A(n_50), .Y(n_877) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_52), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_53), .B(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_54), .A2(n_72), .B1(n_249), .B2(n_535), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_55), .A2(n_75), .B1(n_150), .B2(n_556), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_56), .B(n_199), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_57), .A2(n_154), .B(n_163), .C(n_213), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_58), .A2(n_872), .B1(n_880), .B2(n_881), .Y(n_871) );
INVx1_ASAP7_75t_L g881 ( .A(n_58), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_59), .A2(n_97), .B1(n_533), .B2(n_554), .Y(n_589) );
INVx1_ASAP7_75t_L g146 ( .A(n_60), .Y(n_146) );
AND2x4_ASAP7_75t_L g168 ( .A(n_61), .B(n_169), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_62), .A2(n_63), .B1(n_220), .B2(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_64), .B(n_143), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_65), .B(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_66), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_67), .B(n_220), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_68), .A2(n_105), .B1(n_888), .B2(n_899), .Y(n_104) );
INVx1_ASAP7_75t_L g169 ( .A(n_69), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_70), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_71), .B(n_143), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_73), .B(n_150), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g255 ( .A(n_74), .B(n_200), .C(n_237), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_76), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_77), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_78), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_79), .B(n_165), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_80), .B(n_159), .Y(n_158) );
XNOR2x1_ASAP7_75t_L g131 ( .A(n_81), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g878 ( .A(n_81), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_82), .A2(n_98), .B1(n_163), .B2(n_220), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_83), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_84), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_86), .A2(n_91), .B1(n_194), .B2(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_87), .B(n_165), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g181 ( .A(n_88), .B(n_153), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_89), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_90), .B(n_143), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_92), .Y(n_560) );
INVx1_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_93), .B(n_867), .Y(n_866) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_94), .B(n_165), .Y(n_583) );
INVx1_ASAP7_75t_L g122 ( .A(n_95), .Y(n_122) );
NAND2xp33_ASAP7_75t_L g152 ( .A(n_96), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_99), .B(n_183), .Y(n_203) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_100), .B(n_153), .C(n_176), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_102), .B(n_150), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_103), .B(n_194), .Y(n_197) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_870), .Y(n_105) );
OAI21x1_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_117), .B(n_852), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx12f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_111), .B(n_857), .Y(n_856) );
AND2x2_ASAP7_75t_L g883 ( .A(n_111), .B(n_884), .Y(n_883) );
INVx3_ASAP7_75t_L g886 ( .A(n_111), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_114), .B(n_116), .Y(n_859) );
AND2x6_ASAP7_75t_SL g865 ( .A(n_115), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g892 ( .A(n_116), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B1(n_850), .B2(n_851), .Y(n_117) );
INVx1_ASAP7_75t_L g850 ( .A(n_118), .Y(n_850) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g851 ( .A(n_124), .Y(n_851) );
AOI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_131), .B(n_518), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
INVx8_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx12f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
BUFx8_ASAP7_75t_SL g520 ( .A(n_129), .Y(n_520) );
AND2x2_ASAP7_75t_L g858 ( .A(n_129), .B(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx2_ASAP7_75t_L g896 ( .A(n_130), .Y(n_896) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g873 ( .A(n_133), .Y(n_873) );
NAND4xp75_ASAP7_75t_L g133 ( .A(n_134), .B(n_364), .C(n_437), .D(n_496), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_320), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_290), .Y(n_135) );
OAI221xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_223), .B1(n_262), .B2(n_267), .C(n_271), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI21xp33_ASAP7_75t_SL g271 ( .A1(n_138), .A2(n_272), .B(n_276), .Y(n_271) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_186), .Y(n_138) );
AND2x2_ASAP7_75t_L g317 ( .A(n_139), .B(n_274), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_139), .B(n_328), .Y(n_390) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_170), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g273 ( .A(n_141), .Y(n_273) );
INVx4_ASAP7_75t_L g296 ( .A(n_141), .Y(n_296) );
AND2x2_ASAP7_75t_L g324 ( .A(n_141), .B(n_187), .Y(n_324) );
OR2x2_ASAP7_75t_L g486 ( .A(n_141), .B(n_270), .Y(n_486) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
INVx2_ASAP7_75t_L g627 ( .A(n_143), .Y(n_627) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_SL g166 ( .A(n_144), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_SL g172 ( .A(n_144), .Y(n_172) );
INVx2_ASAP7_75t_L g228 ( .A(n_144), .Y(n_228) );
BUFx3_ASAP7_75t_L g568 ( .A(n_144), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_144), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g576 ( .A(n_144), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_144), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_144), .B(n_629), .Y(n_628) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_157), .B(n_166), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_154), .Y(n_148) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_150), .A2(n_219), .B1(n_220), .B2(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g535 ( .A(n_150), .Y(n_535) );
INVx1_ASAP7_75t_L g554 ( .A(n_150), .Y(n_554) );
INVx4_ASAP7_75t_L g556 ( .A(n_150), .Y(n_556) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_151), .Y(n_153) );
INVx1_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx1_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
INVx2_ASAP7_75t_L g215 ( .A(n_151), .Y(n_215) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
INVx1_ASAP7_75t_L g232 ( .A(n_151), .Y(n_232) );
INVx1_ASAP7_75t_L g285 ( .A(n_151), .Y(n_285) );
INVx2_ASAP7_75t_L g249 ( .A(n_153), .Y(n_249) );
INVx1_ASAP7_75t_L g564 ( .A(n_153), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_154), .A2(n_179), .B(n_181), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_154), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_231), .B(n_233), .Y(n_230) );
BUFx4f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
INVx1_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
BUFx8_ASAP7_75t_L g237 ( .A(n_156), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B1(n_162), .B2(n_164), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_159), .A2(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_165), .A2(n_175), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g259 ( .A(n_165), .Y(n_259) );
INVx3_ASAP7_75t_L g533 ( .A(n_165), .Y(n_533) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_167), .A2(n_174), .B(n_178), .Y(n_173) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_167), .A2(n_191), .B(n_196), .Y(n_190) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_167), .A2(n_230), .B(n_234), .Y(n_229) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_167), .A2(n_242), .B(n_246), .Y(n_241) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_167), .A2(n_253), .B(n_256), .Y(n_252) );
BUFx10_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx10_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
INVx1_ASAP7_75t_L g545 ( .A(n_168), .Y(n_545) );
INVx2_ASAP7_75t_L g299 ( .A(n_170), .Y(n_299) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_170), .Y(n_325) );
INVx1_ASAP7_75t_L g335 ( .A(n_170), .Y(n_335) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g270 ( .A(n_171), .Y(n_270) );
AND2x2_ASAP7_75t_L g426 ( .A(n_171), .B(n_205), .Y(n_426) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_182), .Y(n_171) );
INVx1_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx1_ASAP7_75t_SL g557 ( .A(n_176), .Y(n_557) );
INVx1_ASAP7_75t_L g610 ( .A(n_176), .Y(n_610) );
INVx1_ASAP7_75t_L g565 ( .A(n_180), .Y(n_565) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g189 ( .A(n_184), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_184), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_184), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
INVx2_ASAP7_75t_L g288 ( .A(n_185), .Y(n_288) );
INVx2_ASAP7_75t_L g383 ( .A(n_186), .Y(n_383) );
AND2x2_ASAP7_75t_L g387 ( .A(n_186), .B(n_299), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_186), .B(n_418), .Y(n_516) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_204), .Y(n_186) );
INVx2_ASAP7_75t_L g350 ( .A(n_187), .Y(n_350) );
AND2x2_ASAP7_75t_L g444 ( .A(n_187), .B(n_310), .Y(n_444) );
AND2x2_ASAP7_75t_L g495 ( .A(n_187), .B(n_296), .Y(n_495) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g269 ( .A(n_188), .Y(n_269) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_203), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_241), .B(n_250), .Y(n_240) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_189), .A2(n_241), .B(n_250), .Y(n_266) );
OAI21xp33_ASAP7_75t_SL g275 ( .A1(n_189), .A2(n_190), .B(n_203), .Y(n_275) );
INVx1_ASAP7_75t_L g553 ( .A(n_194), .Y(n_553) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_201), .Y(n_196) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g217 ( .A(n_202), .Y(n_217) );
AND2x2_ASAP7_75t_L g274 ( .A(n_204), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g298 ( .A(n_205), .Y(n_298) );
AOI21x1_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_211), .B(n_222), .Y(n_205) );
NOR2xp67_ASAP7_75t_SL g206 ( .A(n_207), .B(n_209), .Y(n_206) );
INVx2_ASAP7_75t_L g536 ( .A(n_207), .Y(n_536) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_208), .A2(n_210), .A3(n_280), .B(n_286), .Y(n_279) );
NOR2xp33_ASAP7_75t_SL g559 ( .A(n_208), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_208), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g530 ( .A(n_209), .Y(n_530) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AO31x2_ASAP7_75t_L g550 ( .A1(n_210), .A2(n_551), .A3(n_558), .B(n_559), .Y(n_550) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_210), .A2(n_562), .A3(n_568), .B(n_569), .Y(n_561) );
AO31x2_ASAP7_75t_L g623 ( .A1(n_210), .A2(n_624), .A3(n_627), .B(n_628), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_SL g608 ( .A(n_215), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_217), .A2(n_281), .B1(n_283), .B2(n_284), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_217), .A2(n_283), .B1(n_532), .B2(n_534), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_217), .A2(n_283), .B1(n_542), .B2(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_217), .A2(n_283), .B1(n_563), .B2(n_566), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_217), .A2(n_283), .B1(n_625), .B2(n_626), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_239), .Y(n_224) );
INVx2_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
AND2x2_ASAP7_75t_L g427 ( .A(n_225), .B(n_277), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_225), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_225), .B(n_448), .Y(n_457) );
OR2x2_ASAP7_75t_L g480 ( .A(n_225), .B(n_339), .Y(n_480) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_226), .B(n_306), .Y(n_363) );
AND2x2_ASAP7_75t_L g469 ( .A(n_226), .B(n_278), .Y(n_469) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_238), .Y(n_227) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_228), .A2(n_252), .B(n_261), .Y(n_251) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_228), .A2(n_252), .B(n_261), .Y(n_278) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_228), .A2(n_229), .B(n_238), .Y(n_315) );
INVx2_ASAP7_75t_L g244 ( .A(n_232), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .Y(n_234) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_237), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
INVx6_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
O2A1O1Ixp5_ASAP7_75t_L g578 ( .A1(n_237), .A2(n_556), .B(n_579), .C(n_580), .Y(n_578) );
AND2x2_ASAP7_75t_L g356 ( .A(n_239), .B(n_301), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_239), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_239), .B(n_412), .Y(n_420) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_251), .Y(n_239) );
AND2x2_ASAP7_75t_L g332 ( .A(n_240), .B(n_278), .Y(n_332) );
INVx1_ASAP7_75t_L g476 ( .A(n_240), .Y(n_476) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_279), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_251), .B(n_279), .Y(n_397) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g502 ( .A(n_263), .B(n_305), .Y(n_502) );
AND2x2_ASAP7_75t_L g432 ( .A(n_264), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_265), .Y(n_289) );
AND2x2_ASAP7_75t_L g313 ( .A(n_265), .B(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g319 ( .A(n_265), .Y(n_319) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_265), .Y(n_355) );
INVx1_ASAP7_75t_L g380 ( .A(n_265), .Y(n_380) );
AND2x2_ASAP7_75t_L g386 ( .A(n_265), .B(n_278), .Y(n_386) );
INVx1_ASAP7_75t_L g467 ( .A(n_265), .Y(n_467) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_310), .Y(n_309) );
AOI32xp33_ASAP7_75t_SL g441 ( .A1(n_268), .A2(n_333), .A3(n_442), .B1(n_444), .B2(n_445), .Y(n_441) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
OR2x2_ASAP7_75t_L g343 ( .A(n_269), .B(n_299), .Y(n_343) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_270), .Y(n_347) );
INVxp67_ASAP7_75t_L g373 ( .A(n_270), .Y(n_373) );
OR2x2_ASAP7_75t_L g475 ( .A(n_270), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR3x2_ASAP7_75t_L g340 ( .A(n_273), .B(n_341), .C(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g446 ( .A(n_273), .Y(n_446) );
AND2x2_ASAP7_75t_L g374 ( .A(n_274), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g430 ( .A(n_274), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_274), .B(n_325), .Y(n_436) );
BUFx2_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_289), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_277), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_277), .Y(n_509) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g306 ( .A(n_278), .Y(n_306) );
INVx1_ASAP7_75t_L g448 ( .A(n_278), .Y(n_448) );
INVx1_ASAP7_75t_L g307 ( .A(n_279), .Y(n_307) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_279), .Y(n_353) );
OR2x2_ASAP7_75t_L g394 ( .A(n_279), .B(n_315), .Y(n_394) );
AND2x2_ASAP7_75t_L g412 ( .A(n_279), .B(n_315), .Y(n_412) );
AND2x2_ASAP7_75t_L g433 ( .A(n_279), .B(n_303), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_283), .A2(n_552), .B1(n_555), .B2(n_557), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_283), .A2(n_582), .B(n_583), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_283), .A2(n_557), .B1(n_589), .B2(n_590), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_283), .A2(n_607), .B1(n_609), .B2(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g567 ( .A(n_285), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
BUFx2_ASAP7_75t_L g558 ( .A(n_288), .Y(n_558) );
BUFx2_ASAP7_75t_L g501 ( .A(n_289), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_308), .C(n_316), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_300), .Y(n_291) );
INVx3_ASAP7_75t_L g423 ( .A(n_292), .Y(n_423) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g453 ( .A(n_294), .B(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g375 ( .A(n_295), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_295), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g460 ( .A(n_295), .B(n_299), .Y(n_460) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g334 ( .A(n_296), .B(n_335), .Y(n_334) );
NAND2x1_ASAP7_75t_L g349 ( .A(n_296), .B(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g418 ( .A(n_296), .Y(n_418) );
NAND2xp33_ASAP7_75t_R g401 ( .A(n_297), .B(n_324), .Y(n_401) );
AND2x2_ASAP7_75t_L g417 ( .A(n_297), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g483 ( .A(n_297), .Y(n_483) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
INVx1_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
INVx2_ASAP7_75t_L g409 ( .A(n_298), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_299), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g331 ( .A(n_302), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g318 ( .A(n_305), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g489 ( .A(n_305), .B(n_380), .Y(n_489) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g370 ( .A(n_307), .B(n_315), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g337 ( .A(n_313), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g440 ( .A(n_314), .Y(n_440) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g498 ( .A(n_317), .Y(n_498) );
INVx1_ASAP7_75t_L g326 ( .A(n_318), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_319), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g396 ( .A(n_319), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g443 ( .A(n_319), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_319), .B(n_393), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .C(n_344), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g358 ( .A(n_324), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g451 ( .A(n_324), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_336), .B2(n_340), .Y(n_327) );
NAND3x2_ASAP7_75t_L g470 ( .A(n_328), .B(n_471), .C(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_332), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g382 ( .A(n_334), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g454 ( .A(n_334), .Y(n_454) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g506 ( .A(n_338), .B(n_439), .Y(n_506) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
NOR2x1p5_ASAP7_75t_SL g415 ( .A(n_341), .B(n_343), .Y(n_415) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g359 ( .A(n_342), .Y(n_359) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_342), .Y(n_461) );
OAI22xp33_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_351), .B1(n_357), .B2(n_360), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g504 ( .A(n_347), .B(n_451), .Y(n_504) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OR2x6_ASAP7_75t_L g424 ( .A(n_349), .B(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_356), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g406 ( .A(n_353), .Y(n_406) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_358), .A2(n_474), .B1(n_479), .B2(n_481), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_358), .A2(n_452), .B1(n_509), .B2(n_510), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_358), .B(n_506), .Y(n_513) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_365), .B(n_398), .Y(n_364) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_376), .C(n_388), .Y(n_365) );
AO21x1_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g468 ( .A(n_367), .Y(n_468) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
AOI32xp33_ASAP7_75t_L g488 ( .A1(n_372), .A2(n_489), .A3(n_490), .B1(n_491), .B2(n_493), .Y(n_488) );
BUFx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g471 ( .A(n_375), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_384), .B2(n_387), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g404 ( .A(n_380), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_380), .B(n_412), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_381), .A2(n_389), .B1(n_391), .B2(n_395), .Y(n_388) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g485 ( .A(n_383), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI322xp33_ASAP7_75t_L g497 ( .A1(n_385), .A2(n_478), .A3(n_498), .B1(n_499), .B2(n_503), .C1(n_504), .C2(n_505), .Y(n_497) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g517 ( .A(n_386), .B(n_406), .Y(n_517) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g478 ( .A(n_394), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g435 ( .A(n_397), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_421), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B(n_407), .C(n_416), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_413), .B2(n_414), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_412), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_412), .B(n_448), .Y(n_511) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_427), .B(n_428), .Y(n_421) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NOR2x1_ASAP7_75t_SL g450 ( .A(n_425), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g487 ( .A(n_427), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_434), .B2(n_436), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NOR3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_462), .C(n_484), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B(n_449), .C(n_458), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g456 ( .A(n_443), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_444), .B(n_446), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_452), .B(n_455), .Y(n_449) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVxp67_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_470), .B(n_473), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .C(n_469), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OAI21xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_487), .B(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .C(n_512), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
AND3x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_747), .C(n_825), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_690), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_637), .C(n_660), .Y(n_523) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_571), .B1(n_593), .B2(n_602), .C(n_613), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_548), .Y(n_525) );
AND2x4_ASAP7_75t_L g727 ( .A(n_526), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
INVx2_ASAP7_75t_L g686 ( .A(n_528), .Y(n_686) );
INVx1_ASAP7_75t_L g713 ( .A(n_528), .Y(n_713) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g596 ( .A(n_529), .Y(n_596) );
AND2x4_ASAP7_75t_L g664 ( .A(n_529), .B(n_597), .Y(n_664) );
AO31x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .A3(n_536), .B(n_537), .Y(n_529) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_530), .A2(n_558), .A3(n_588), .B(n_591), .Y(n_587) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_536), .A2(n_541), .A3(n_544), .B(n_546), .Y(n_540) );
INVx1_ASAP7_75t_L g746 ( .A(n_539), .Y(n_746) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g597 ( .A(n_540), .Y(n_597) );
AND2x4_ASAP7_75t_L g635 ( .A(n_540), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g655 ( .A(n_540), .B(n_561), .Y(n_655) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_540), .Y(n_707) );
INVx1_ASAP7_75t_L g800 ( .A(n_540), .Y(n_800) );
AND2x2_ASAP7_75t_L g846 ( .A(n_540), .B(n_550), .Y(n_846) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_544), .A2(n_568), .A3(n_606), .B(n_611), .Y(n_605) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g584 ( .A(n_545), .Y(n_584) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_549), .B(n_712), .Y(n_711) );
NAND2x1_ASAP7_75t_L g716 ( .A(n_549), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g840 ( .A(n_549), .B(n_738), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_549), .B(n_794), .Y(n_844) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_561), .Y(n_549) );
INVx4_ASAP7_75t_SL g599 ( .A(n_550), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_550), .B(n_601), .Y(n_648) );
BUFx2_ASAP7_75t_L g732 ( .A(n_550), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_550), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
INVx2_ASAP7_75t_L g636 ( .A(n_561), .Y(n_636) );
AND2x2_ASAP7_75t_L g638 ( .A(n_561), .B(n_596), .Y(n_638) );
INVx1_ASAP7_75t_L g663 ( .A(n_561), .Y(n_663) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_561), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_561), .B(n_746), .Y(n_777) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g821 ( .A(n_573), .B(n_822), .Y(n_821) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_586), .Y(n_573) );
AND2x4_ASAP7_75t_L g617 ( .A(n_574), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g678 ( .A(n_574), .B(n_622), .Y(n_678) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g764 ( .A(n_575), .Y(n_764) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_585), .Y(n_575) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_576), .A2(n_577), .B(n_585), .Y(n_651) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_584), .Y(n_577) );
AND2x4_ASAP7_75t_L g676 ( .A(n_586), .B(n_605), .Y(n_676) );
INVx3_ASAP7_75t_L g699 ( .A(n_586), .Y(n_699) );
INVx2_ASAP7_75t_L g720 ( .A(n_586), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_586), .B(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_586), .B(n_621), .Y(n_814) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g604 ( .A(n_587), .B(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g616 ( .A(n_587), .Y(n_616) );
AND2x2_ASAP7_75t_L g693 ( .A(n_587), .B(n_618), .Y(n_693) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx3_ASAP7_75t_L g671 ( .A(n_596), .Y(n_671) );
AND2x2_ASAP7_75t_L g706 ( .A(n_596), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g775 ( .A(n_596), .B(n_599), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_597), .B(n_599), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_598), .B(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g634 ( .A(n_599), .Y(n_634) );
AND2x2_ASAP7_75t_L g662 ( .A(n_599), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g680 ( .A(n_599), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g722 ( .A(n_599), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_599), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g783 ( .A(n_599), .Y(n_783) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_604), .B(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_SL g657 ( .A(n_604), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g736 ( .A(n_604), .B(n_620), .Y(n_736) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_604), .Y(n_771) );
INVx2_ASAP7_75t_L g788 ( .A(n_604), .Y(n_788) );
INVx2_ASAP7_75t_L g618 ( .A(n_605), .Y(n_618) );
OR2x2_ASAP7_75t_L g668 ( .A(n_605), .B(n_659), .Y(n_668) );
INVx1_ASAP7_75t_L g689 ( .A(n_605), .Y(n_689) );
BUFx2_ASAP7_75t_L g704 ( .A(n_605), .Y(n_704) );
OR2x2_ASAP7_75t_L g773 ( .A(n_605), .B(n_623), .Y(n_773) );
AOI21xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_619), .B(n_631), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g739 ( .A1(n_614), .A2(n_695), .B(n_740), .C(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g639 ( .A(n_615), .B(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_615), .A2(n_673), .B1(n_839), .B2(n_840), .Y(n_838) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
AND2x4_ASAP7_75t_L g758 ( .A(n_617), .B(n_667), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_617), .B(n_813), .Y(n_812) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_630), .Y(n_619) );
INVx1_ASAP7_75t_L g640 ( .A(n_620), .Y(n_640) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_L g658 ( .A(n_621), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_622), .B(n_651), .Y(n_701) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g650 ( .A(n_623), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g667 ( .A(n_623), .Y(n_667) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_623), .Y(n_742) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
AND2x2_ASAP7_75t_L g653 ( .A(n_633), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_634), .B(n_713), .Y(n_752) );
INVx2_ASAP7_75t_L g644 ( .A(n_635), .Y(n_644) );
AND2x2_ASAP7_75t_L g721 ( .A(n_635), .B(n_722), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_635), .B(n_685), .Y(n_766) );
AND2x2_ASAP7_75t_L g803 ( .A(n_635), .B(n_775), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_641), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_649), .B1(n_652), .B2(n_656), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g847 ( .A(n_644), .Y(n_847) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g687 ( .A(n_650), .Y(n_687) );
AND2x2_ASAP7_75t_L g714 ( .A(n_650), .B(n_699), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_650), .B(n_693), .Y(n_784) );
AND2x4_ASAP7_75t_L g830 ( .A(n_650), .B(n_676), .Y(n_830) );
INVx1_ASAP7_75t_L g659 ( .A(n_651), .Y(n_659) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g836 ( .A(n_654), .B(n_732), .Y(n_836) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g769 ( .A(n_655), .B(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_L g797 ( .A(n_655), .B(n_671), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_656), .B(n_829), .Y(n_828) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g778 ( .A(n_658), .B(n_779), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_665), .B1(n_669), .B2(n_673), .C(n_679), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g695 ( .A(n_662), .Y(n_695) );
AND2x2_ASAP7_75t_L g819 ( .A(n_662), .B(n_685), .Y(n_819) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_663), .Y(n_683) );
INVx3_ASAP7_75t_L g681 ( .A(n_664), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_664), .B(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g753 ( .A(n_664), .B(n_754), .Y(n_753) );
NOR2xp67_ASAP7_75t_SL g665 ( .A(n_666), .B(n_668), .Y(n_665) );
AND2x2_ASAP7_75t_L g692 ( .A(n_666), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_666), .B(n_699), .Y(n_761) );
AOI322xp5_ASAP7_75t_L g767 ( .A1(n_666), .A2(n_753), .A3(n_768), .B1(n_771), .B2(n_772), .C1(n_774), .C2(n_778), .Y(n_767) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g709 ( .A(n_667), .B(n_676), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_668), .B(n_720), .Y(n_719) );
NOR2x1_ASAP7_75t_L g817 ( .A(n_668), .B(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_669), .A2(n_811), .B1(n_815), .B2(n_819), .Y(n_810) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx4_ASAP7_75t_L g794 ( .A(n_671), .Y(n_794) );
OR2x2_ASAP7_75t_L g824 ( .A(n_671), .B(n_799), .Y(n_824) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g837 ( .A(n_676), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_677), .B(n_703), .Y(n_724) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI211x1_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B(n_687), .C(n_688), .Y(n_679) );
INVx2_ASAP7_75t_L g717 ( .A(n_681), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g744 ( .A(n_685), .Y(n_744) );
NAND2x1_ASAP7_75t_L g835 ( .A(n_685), .B(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g741 ( .A(n_686), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g806 ( .A(n_688), .Y(n_806) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_708), .C(n_723), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_696), .C(n_706), .Y(n_691) );
INVx1_ASAP7_75t_L g705 ( .A(n_692), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_693), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g763 ( .A(n_693), .B(n_764), .Y(n_763) );
NAND2xp33_ASAP7_75t_L g786 ( .A(n_693), .B(n_734), .Y(n_786) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_705), .Y(n_696) );
INVx1_ASAP7_75t_L g832 ( .A(n_697), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g779 ( .A(n_699), .Y(n_779) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g734 ( .A(n_701), .Y(n_734) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_701), .Y(n_809) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g738 ( .A(n_707), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_714), .B2(n_715), .C(n_718), .Y(n_708) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g770 ( .A(n_713), .Y(n_770) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g756 ( .A(n_720), .Y(n_756) );
NOR2x1p5_ASAP7_75t_L g772 ( .A(n_720), .B(n_773), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_721), .A2(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g728 ( .A(n_722), .Y(n_728) );
AOI211xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B(n_729), .C(n_739), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_733), .B1(n_735), .B2(n_737), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g818 ( .A(n_742), .Y(n_818) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_780), .C(n_801), .Y(n_747) );
NAND3xp33_ASAP7_75t_SL g748 ( .A(n_749), .B(n_759), .C(n_767), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B(n_755), .Y(n_749) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
AND2x2_ASAP7_75t_L g849 ( .A(n_756), .B(n_817), .Y(n_849) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g795 ( .A1(n_758), .A2(n_796), .B(n_798), .Y(n_795) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
OR2x2_ASAP7_75t_L g787 ( .A(n_764), .B(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g822 ( .A(n_773), .Y(n_822) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_776), .Y(n_839) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g782 ( .A(n_777), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g792 ( .A(n_777), .Y(n_792) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_784), .B1(n_785), .B2(n_789), .C(n_795), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_781), .A2(n_827), .B(n_831), .Y(n_826) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI32xp33_ASAP7_75t_L g820 ( .A1(n_783), .A2(n_794), .A3(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
AND2x2_ASAP7_75t_SL g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_796), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI211xp5_ASAP7_75t_SL g801 ( .A1(n_802), .A2(n_804), .B(n_810), .C(n_820), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_833), .C(n_841), .Y(n_825) );
INVxp33_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI21xp33_ASAP7_75t_SL g833 ( .A1(n_834), .A2(n_837), .B(n_838), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_845), .B(n_848), .Y(n_841) );
INVxp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NOR2xp33_ASAP7_75t_SL g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
BUFx10_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVxp67_ASAP7_75t_SL g887 ( .A(n_860), .Y(n_887) );
NOR2xp67_ASAP7_75t_SL g860 ( .A(n_861), .B(n_869), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
INVx4_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx12f_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx4_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx5_ASAP7_75t_L g884 ( .A(n_865), .Y(n_884) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_868), .Y(n_894) );
OAI22x1_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_882), .B1(n_885), .B2(n_887), .Y(n_870) );
INVx2_ASAP7_75t_L g880 ( .A(n_872), .Y(n_880) );
XNOR2x1_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_883), .Y(n_882) );
BUFx8_ASAP7_75t_SL g885 ( .A(n_886), .Y(n_885) );
BUFx12f_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_889), .Y(n_899) );
INVx6_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
NAND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_892), .Y(n_891) );
NOR2x1p5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
endmodule