module fake_jpeg_1586_n_388 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_8),
.B(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_47),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_20),
.B(n_0),
.CON(n_52),
.SN(n_52)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_85),
.B(n_0),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_59),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_72),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_69),
.B(n_80),
.Y(n_121)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_76),
.B(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

CKINVDCx9p33_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_84),
.B1(n_18),
.B2(n_41),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_1),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_70),
.B1(n_51),
.B2(n_64),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_18),
.B1(n_41),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_90),
.A2(n_96),
.B1(n_114),
.B2(n_122),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_93),
.A2(n_95),
.B1(n_103),
.B2(n_79),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_16),
.C(n_17),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_129),
.C(n_76),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_27),
.B1(n_41),
.B2(n_39),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_107),
.B1(n_109),
.B2(n_118),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_26),
.B1(n_39),
.B2(n_35),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g177 ( 
.A1(n_99),
.A2(n_11),
.B1(n_7),
.B2(n_9),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_16),
.B1(n_35),
.B2(n_34),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_105),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_16),
.B1(n_34),
.B2(n_33),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_32),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_112),
.B(n_127),
.CON(n_158),
.SN(n_158)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_22),
.B1(n_42),
.B2(n_16),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_71),
.A2(n_16),
.B1(n_22),
.B2(n_42),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_126),
.B1(n_94),
.B2(n_127),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_16),
.B1(n_42),
.B2(n_3),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_57),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

FAx1_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_15),
.CI(n_14),
.CON(n_127),
.SN(n_127)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_65),
.B(n_1),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_4),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_140),
.A2(n_176),
.B1(n_179),
.B2(n_115),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_75),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_142),
.B(n_153),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_174),
.B1(n_178),
.B2(n_105),
.Y(n_188)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_85),
.B1(n_77),
.B2(n_83),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_148),
.A2(n_150),
.B1(n_154),
.B2(n_152),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_156),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_80),
.B1(n_81),
.B2(n_78),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_118),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_14),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_154),
.B(n_157),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_91),
.A3(n_132),
.B1(n_131),
.B2(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_159),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_13),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_12),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_84),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_84),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_167),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_171),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_99),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_5),
.C(n_6),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_177),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_89),
.B(n_6),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_97),
.B(n_7),
.Y(n_178)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_135),
.Y(n_198)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_183),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_92),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_200),
.B(n_152),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_146),
.B1(n_141),
.B2(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_187),
.A2(n_207),
.B1(n_140),
.B2(n_113),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_188),
.B(n_177),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_91),
.B1(n_134),
.B2(n_106),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_202),
.B1(n_180),
.B2(n_147),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_134),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_106),
.B1(n_107),
.B2(n_125),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_212),
.B1(n_196),
.B2(n_198),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_141),
.A2(n_135),
.B1(n_125),
.B2(n_115),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_124),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_130),
.B1(n_128),
.B2(n_116),
.Y(n_212)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_205),
.B(n_197),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_219),
.A2(n_207),
.B(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_138),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_139),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_228),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_174),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_227),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_168),
.C(n_162),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_209),
.C(n_189),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_178),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_231),
.B(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_160),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_158),
.B(n_177),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_239),
.B(n_189),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_158),
.B(n_140),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_185),
.A2(n_152),
.B(n_140),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_246),
.B(n_196),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_248),
.B1(n_249),
.B2(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_185),
.B(n_177),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_203),
.A2(n_128),
.B1(n_130),
.B2(n_102),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_263),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_226),
.Y(n_281)
);

AO22x1_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_196),
.B1(n_200),
.B2(n_186),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_271),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_261),
.B(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_184),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_269),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_265),
.C(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_195),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_196),
.B1(n_181),
.B2(n_195),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_275),
.B1(n_221),
.B2(n_254),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_276),
.B1(n_249),
.B2(n_237),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_233),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_230),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_181),
.B1(n_204),
.B2(n_218),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_219),
.A2(n_145),
.B1(n_102),
.B2(n_116),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_258),
.A2(n_239),
.B(n_236),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_282),
.B(n_250),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_296),
.C(n_259),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_238),
.B(n_236),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_254),
.B1(n_276),
.B2(n_259),
.Y(n_301)
);

NOR4xp25_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_228),
.C(n_231),
.D(n_241),
.Y(n_285)
);

OA21x2_ASAP7_75t_SL g316 ( 
.A1(n_285),
.A2(n_294),
.B(n_283),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_239),
.B1(n_246),
.B2(n_220),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_298),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_224),
.B1(n_226),
.B2(n_237),
.Y(n_289)
);

BUFx12f_ASAP7_75t_SL g290 ( 
.A(n_252),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_292),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_257),
.A2(n_251),
.B(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_245),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_245),
.C(n_235),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_297),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_225),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_240),
.B1(n_244),
.B2(n_210),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_270),
.B1(n_263),
.B2(n_260),
.Y(n_315)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_301),
.A2(n_305),
.B1(n_310),
.B2(n_312),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_311),
.C(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_256),
.B1(n_277),
.B2(n_261),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_293),
.B1(n_288),
.B2(n_282),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_315),
.B1(n_319),
.B2(n_278),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_256),
.B1(n_277),
.B2(n_265),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_291),
.C(n_296),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_257),
.B1(n_270),
.B2(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_292),
.C(n_279),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_279),
.C(n_278),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_257),
.B1(n_260),
.B2(n_274),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_290),
.B(n_295),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_332),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_303),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_329),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_325),
.B(n_316),
.Y(n_343)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_302),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_327),
.A2(n_305),
.B1(n_319),
.B2(n_312),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_286),
.C(n_283),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_335),
.C(n_336),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_234),
.B(n_208),
.Y(n_347)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

BUFx12_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

NAND4xp25_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_337),
.C(n_309),
.D(n_242),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_286),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_208),
.C(n_218),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_341),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_327),
.A2(n_301),
.B1(n_309),
.B2(n_314),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_343),
.B(n_345),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_322),
.A2(n_324),
.B1(n_334),
.B2(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_300),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_318),
.B1(n_320),
.B2(n_247),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_329),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_347),
.A2(n_333),
.B(n_234),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_335),
.A2(n_210),
.B1(n_204),
.B2(n_234),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_349),
.B(n_351),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_328),
.C(n_323),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_321),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_354),
.Y(n_368)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_350),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_336),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_355),
.B(n_345),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_346),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_357),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_347),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_328),
.B(n_333),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_SL g363 ( 
.A(n_362),
.B(n_350),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_169),
.B(n_144),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_359),
.B(n_354),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_366),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_361),
.A2(n_339),
.B1(n_341),
.B2(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_172),
.C(n_182),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_340),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_371),
.A2(n_213),
.B(n_182),
.Y(n_374)
);

AOI321xp33_ASAP7_75t_L g373 ( 
.A1(n_368),
.A2(n_356),
.A3(n_361),
.B1(n_352),
.B2(n_213),
.C(n_183),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_373),
.A2(n_364),
.B(n_214),
.C(n_194),
.Y(n_379)
);

OAI31xp33_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_378),
.A3(n_214),
.B(n_163),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_367),
.A2(n_217),
.B(n_215),
.C(n_194),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_163),
.B(n_101),
.C(n_364),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_379),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_380),
.A2(n_382),
.B1(n_163),
.B2(n_108),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_385),
.C(n_9),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_372),
.A3(n_376),
.B1(n_172),
.B2(n_124),
.C1(n_108),
.C2(n_7),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_386),
.B(n_383),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_9),
.Y(n_388)
);


endmodule