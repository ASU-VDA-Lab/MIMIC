module fake_jpeg_19162_n_376 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_376);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_376;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_1),
.B(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_69),
.Y(n_85)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_48),
.B(n_53),
.Y(n_115)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_49),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_16),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_56),
.B(n_58),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_65),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_62),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_132)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_3),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_18),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_77),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_4),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_23),
.C(n_26),
.Y(n_100)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_4),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_44),
.B1(n_21),
.B2(n_35),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_88),
.B1(n_94),
.B2(n_117),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_93),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_22),
.B1(n_36),
.B2(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_96),
.B(n_111),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_24),
.B(n_29),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_38),
.C(n_33),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_108),
.B1(n_119),
.B2(n_62),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_96),
.B1(n_103),
.B2(n_99),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_123),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_81),
.B1(n_67),
.B2(n_54),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_23),
.B1(n_18),
.B2(n_38),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_48),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_7),
.Y(n_170)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_133),
.B1(n_90),
.B2(n_105),
.Y(n_187)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_138),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_155),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_75),
.B1(n_77),
.B2(n_71),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_172),
.B1(n_126),
.B2(n_92),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_84),
.Y(n_183)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_55),
.C(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_99),
.A2(n_38),
.B1(n_33),
.B2(n_9),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_85),
.B(n_38),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_61),
.B(n_64),
.C(n_82),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_158),
.A2(n_164),
.B1(n_130),
.B2(n_91),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_80),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_176),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_72),
.B1(n_70),
.B2(n_68),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_170),
.Y(n_202)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

CKINVDCx6p67_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_10),
.C(n_11),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_122),
.C(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_88),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_183),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_90),
.B1(n_133),
.B2(n_105),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_187),
.B1(n_192),
.B2(n_198),
.Y(n_230)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_87),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_130),
.B1(n_118),
.B2(n_86),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_121),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_121),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_141),
.A2(n_131),
.B(n_11),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_10),
.B(n_12),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_207),
.B1(n_210),
.B2(n_156),
.Y(n_228)
);

AND2x4_ASAP7_75t_SL g203 ( 
.A(n_158),
.B(n_122),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_194),
.B1(n_200),
.B2(n_191),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_134),
.A2(n_157),
.B1(n_165),
.B2(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_149),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_101),
.B1(n_86),
.B2(n_13),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_138),
.B1(n_159),
.B2(n_145),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_153),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_138),
.B1(n_152),
.B2(n_150),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_143),
.A2(n_101),
.B1(n_12),
.B2(n_13),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_222),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_144),
.B1(n_161),
.B2(n_169),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_184),
.B(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_160),
.B1(n_135),
.B2(n_174),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_171),
.B1(n_166),
.B2(n_142),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_201),
.B1(n_196),
.B2(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_149),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_245),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_178),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_213),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_247),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_147),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_221),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_198),
.B1(n_192),
.B2(n_194),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_271),
.B1(n_230),
.B2(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_194),
.C(n_179),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_225),
.C(n_239),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_265),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_248),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_188),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_267),
.B(n_220),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_196),
.B(n_223),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_245),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_202),
.B1(n_181),
.B2(n_210),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_217),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_274),
.B(n_283),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_284),
.B(n_295),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_294),
.B(n_296),
.C(n_261),
.Y(n_297)
);

AOI221xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_219),
.B1(n_232),
.B2(n_221),
.C(n_215),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_230),
.B1(n_237),
.B2(n_235),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_202),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_225),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_225),
.B(n_246),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_292),
.C(n_252),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_215),
.B1(n_242),
.B2(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_254),
.B1(n_271),
.B2(n_266),
.Y(n_306)
);

OAI22x1_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_234),
.B1(n_222),
.B2(n_244),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_256),
.B1(n_273),
.B2(n_216),
.Y(n_313)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_266),
.C(n_260),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_247),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_262),
.A2(n_224),
.B(n_202),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_254),
.A2(n_243),
.B(n_233),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_296),
.B(n_290),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_309),
.C(n_283),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_303),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_259),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_264),
.B1(n_260),
.B2(n_259),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_311),
.B1(n_313),
.B2(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_272),
.C(n_262),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_284),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_272),
.A3(n_263),
.B1(n_273),
.B2(n_269),
.C1(n_250),
.C2(n_229),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_293),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_310),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_317),
.A2(n_324),
.B(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_285),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_321),
.A2(n_323),
.B1(n_298),
.B2(n_319),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_276),
.B1(n_278),
.B2(n_287),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_315),
.B1(n_307),
.B2(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_280),
.B1(n_282),
.B2(n_277),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_280),
.B(n_275),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_294),
.B(n_288),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_325),
.A2(n_329),
.B(n_307),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_286),
.C(n_283),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_311),
.A2(n_291),
.B(n_263),
.C(n_295),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_304),
.A2(n_279),
.B(n_292),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_189),
.C(n_206),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_331),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_343),
.B1(n_328),
.B2(n_314),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_325),
.A2(n_309),
.B1(n_300),
.B2(n_301),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_335),
.A2(n_322),
.B(n_142),
.Y(n_353)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_337),
.A2(n_317),
.B(n_324),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_316),
.C(n_326),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_303),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_341),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_310),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_308),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_323),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_258),
.B1(n_314),
.B2(n_181),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_352),
.C(n_354),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_347),
.A2(n_338),
.B(n_344),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_351),
.Y(n_363)
);

AOI211xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_321),
.B(n_319),
.C(n_329),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g355 ( 
.A1(n_350),
.A2(n_335),
.B(n_338),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_318),
.C(n_331),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_353),
.A2(n_181),
.B1(n_206),
.B2(n_147),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_258),
.B1(n_181),
.B2(n_238),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_355),
.A2(n_360),
.B(n_12),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_SL g356 ( 
.A(n_347),
.B(n_334),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_357),
.B(n_362),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_339),
.C(n_340),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_346),
.C(n_353),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_349),
.A2(n_342),
.B(n_341),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_352),
.B(n_114),
.Y(n_361)
);

AOI211xp5_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_12),
.B(n_13),
.C(n_109),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_351),
.C(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_238),
.C(n_114),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_367),
.A2(n_369),
.B(n_357),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_368),
.A2(n_13),
.B1(n_112),
.B2(n_365),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_373),
.C(n_372),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_371),
.Y(n_376)
);


endmodule