module real_jpeg_1678_n_29 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_156, n_24, n_165, n_6, n_159, n_28, n_161, n_162, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_155, n_29);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_156;
input n_24;
input n_165;
input n_6;
input n_159;
input n_28;
input n_161;
input n_162;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_74;
wire n_41;
wire n_32;
wire n_80;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_2),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_3),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_4),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_6),
.B(n_51),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_77),
.B(n_81),
.Y(n_76)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_8),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_144),
.B2(n_147),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_9),
.B(n_33),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.C(n_95),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_12),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_17),
.A2(n_68),
.B1(n_101),
.B2(n_104),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_19),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_72),
.C(n_87),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_75),
.B2(n_86),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_28),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_150),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_41),
.B(n_143),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_37),
.B(n_136),
.Y(n_135)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_37),
.Y(n_149)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_74),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_40),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_40),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_139),
.C(n_140),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_138),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_44),
.B(n_47),
.Y(n_138)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B(n_54),
.C(n_137),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_53),
.B(n_153),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_133),
.C(n_134),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_132),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_142),
.Y(n_141)
);

OAI221xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_107),
.C(n_122),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_97),
.C(n_98),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_90),
.C(n_91),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.C(n_85),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_123),
.A3(n_124),
.B1(n_127),
.B2(n_128),
.C1(n_131),
.C2(n_165),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.C(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_155),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_156),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_157),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_158),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_159),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_160),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_161),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_162),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_163),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_164),
.Y(n_121)
);


endmodule