module fake_jpeg_27943_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_45),
.B1(n_23),
.B2(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_61),
.B1(n_69),
.B2(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_23),
.B1(n_15),
.B2(n_24),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_15),
.B1(n_24),
.B2(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_85),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_15),
.CI(n_32),
.CON(n_80),
.SN(n_80)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_104),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_65),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_32),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_63),
.B(n_27),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_26),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_59),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_64),
.B1(n_71),
.B2(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_120),
.B1(n_96),
.B2(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_121),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_74),
.B1(n_67),
.B2(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_98),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_75),
.B(n_62),
.C(n_63),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_116),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_1),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_121),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.C(n_95),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_10),
.C(n_5),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_81),
.C(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_103),
.B1(n_80),
.B2(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_97),
.B1(n_91),
.B2(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_96),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_7),
.B(n_8),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_125),
.B(n_126),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_8),
.C(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_123),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_116),
.B(n_113),
.C(n_124),
.D(n_105),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_128),
.B(n_141),
.C(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_157),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_126),
.B(n_114),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_142),
.B1(n_143),
.B2(n_128),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_111),
.A3(n_114),
.B1(n_118),
.B2(n_119),
.C1(n_123),
.C2(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_162),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_133),
.C(n_138),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_132),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_163),
.CI(n_164),
.CON(n_181),
.SN(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_149),
.B1(n_161),
.B2(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_150),
.A3(n_148),
.B1(n_159),
.B2(n_144),
.C1(n_161),
.C2(n_156),
.Y(n_178)
);

AOI22x1_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_134),
.B1(n_139),
.B2(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_172),
.B1(n_166),
.B2(n_169),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_149),
.B1(n_157),
.B2(n_134),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_180),
.B(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_156),
.B1(n_111),
.B2(n_118),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_188),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_171),
.C(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_180),
.B(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_175),
.C(n_182),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_194),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_192),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_190),
.C(n_195),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_195),
.Y(n_202)
);


endmodule