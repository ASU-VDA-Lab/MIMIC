module real_jpeg_33413_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_675;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_0),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_1),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_3),
.A2(n_215),
.B1(n_236),
.B2(n_242),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_3),
.A2(n_215),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_3),
.A2(n_215),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_4),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_111),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_4),
.A2(n_111),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g654 ( 
.A1(n_4),
.A2(n_111),
.B1(n_622),
.B2(n_655),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_5),
.A2(n_188),
.B1(n_189),
.B2(n_193),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_5),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_5),
.A2(n_108),
.B1(n_188),
.B2(n_345),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_5),
.A2(n_188),
.B1(n_440),
.B2(n_443),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_5),
.A2(n_188),
.B1(n_516),
.B2(n_520),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_6),
.A2(n_169),
.B1(n_286),
.B2(n_291),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_6),
.A2(n_169),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_6),
.A2(n_169),
.B1(n_468),
.B2(n_472),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_7),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_7),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_7),
.B(n_174),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_7),
.A2(n_363),
.B1(n_501),
.B2(n_504),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g590 ( 
.A1(n_7),
.A2(n_145),
.B(n_525),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_11),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_11),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_11),
.A2(n_276),
.B1(n_376),
.B2(n_380),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_11),
.A2(n_276),
.B1(n_492),
.B2(n_496),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_11),
.A2(n_276),
.B1(n_574),
.B2(n_577),
.Y(n_573)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_12),
.Y(n_545)
);

OAI221xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B1(n_640),
.B2(n_675),
.C(n_679),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_13),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_14),
.A2(n_37),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_14),
.A2(n_37),
.B1(n_502),
.B2(n_627),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_16),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_16),
.A2(n_78),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_16),
.A2(n_78),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_16),
.A2(n_78),
.B1(n_616),
.B2(n_622),
.Y(n_615)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_17),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_18),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_18),
.A2(n_59),
.B1(n_67),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_18),
.A2(n_67),
.B1(n_662),
.B2(n_663),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_20),
.B(n_680),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_606),
.B(n_638),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_423),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_355),
.B(n_419),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_300),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_25),
.A2(n_420),
.B(n_421),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_25),
.B(n_300),
.C(n_425),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_248),
.B(n_251),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_224),
.Y(n_26)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_27),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_27),
.A2(n_224),
.B1(n_249),
.B2(n_250),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_118),
.B1(n_119),
.B2(n_223),
.Y(n_27)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_28),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_28),
.B(n_118),
.C(n_249),
.Y(n_608)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_117),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_71),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_30),
.B(n_71),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_40),
.B1(n_62),
.B2(n_70),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_32),
.A2(n_41),
.B1(n_128),
.B2(n_129),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_36),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_39),
.Y(n_125)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g366 ( 
.A1(n_40),
.A2(n_70),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_40),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_40),
.A2(n_488),
.B1(n_489),
.B2(n_490),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_40),
.B(n_556),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g631 ( 
.A1(n_40),
.A2(n_62),
.B(n_70),
.Y(n_631)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_41),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_41),
.A2(n_122),
.B1(n_128),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_41),
.A2(n_491),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g540 ( 
.A(n_43),
.Y(n_540)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_45),
.Y(n_453)
);

OAI22x1_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_47),
.Y(n_551)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_53),
.Y(n_330)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_54),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_55),
.Y(n_263)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_60),
.Y(n_524)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_61),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_61),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_64),
.Y(n_372)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_65),
.Y(n_497)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_66),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_66),
.Y(n_464)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_70),
.B(n_368),
.Y(n_447)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_70),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_84),
.B1(n_107),
.B2(n_115),
.Y(n_71)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_72),
.A2(n_84),
.B1(n_211),
.B2(n_220),
.Y(n_210)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_76),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_83),
.Y(n_315)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_83),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_84),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_84),
.A2(n_115),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_84),
.B(n_285),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_84),
.A2(n_107),
.B1(n_115),
.B2(n_626),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_84),
.B(n_626),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_90),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_96),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g446 ( 
.A(n_97),
.Y(n_446)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_105),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_110),
.Y(n_379)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_110),
.Y(n_504)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_116),
.A2(n_283),
.B1(n_284),
.B2(n_295),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_116),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_R g528 ( 
.A(n_116),
.B(n_363),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_116),
.A2(n_660),
.B(n_665),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_117),
.A2(n_611),
.B1(n_633),
.B2(n_634),
.Y(n_610)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_117),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_160),
.B(n_221),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_120),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_135),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_121),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_128),
.Y(n_488)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2x2_ASAP7_75t_L g351 ( 
.A(n_135),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_145),
.B1(n_151),
.B2(n_155),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_136),
.A2(n_145),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_138),
.Y(n_537)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_139),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_139),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_139),
.Y(n_549)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_145),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_145),
.A2(n_328),
.B1(n_389),
.B2(n_394),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_145),
.A2(n_515),
.B(n_525),
.Y(n_514)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_146),
.A2(n_261),
.B1(n_327),
.B2(n_334),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_146),
.B(n_467),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_146),
.A2(n_568),
.B1(n_571),
.B2(n_572),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_149),
.Y(n_395)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g527 ( 
.A(n_150),
.Y(n_527)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_153),
.Y(n_391)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_R g259 ( 
.A(n_158),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_159),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_209),
.Y(n_160)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_161),
.A2(n_209),
.B1(n_210),
.B2(n_222),
.Y(n_254)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_186),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_162),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_168),
.Y(n_623)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

AO22x1_ASAP7_75t_SL g274 ( 
.A1(n_174),
.A2(n_187),
.B1(n_196),
.B2(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_174),
.B(n_275),
.Y(n_341)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_181),
.B2(n_183),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_185),
.Y(n_294)
);

NAND2x1_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_192),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_192),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_198),
.B1(n_202),
.B2(n_205),
.Y(n_197)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_196),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_196),
.Y(n_614)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_205),
.Y(n_321)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_208),
.Y(n_621)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_220),
.B(n_285),
.Y(n_349)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_225),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_226),
.A2(n_231),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_230),
.Y(n_570)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_233),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_246),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_245),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_235),
.A2(n_245),
.B1(n_613),
.B2(n_615),
.Y(n_612)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_239),
.Y(n_657)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_242),
.Y(n_362)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_245),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_247),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_251),
.B(n_422),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_296),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_253),
.B(n_297),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_255),
.B(n_354),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_274),
.C(n_282),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_R g302 ( 
.A1(n_256),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_268),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_257),
.B(n_268),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_266),
.Y(n_474)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_267),
.Y(n_519)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_271),
.Y(n_442)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_282),
.Y(n_303)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_289),
.Y(n_462)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_290),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_290),
.Y(n_629)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_344),
.B(n_349),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_295),
.A2(n_349),
.B(n_500),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_298),
.A2(n_636),
.B(n_637),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_353),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_301),
.B(n_353),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.C(n_350),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_303),
.A2(n_304),
.B1(n_351),
.B2(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_305),
.B(n_307),
.Y(n_416)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_339),
.C(n_342),
.Y(n_307)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_326),
.Y(n_308)
);

XOR2x2_ASAP7_75t_L g382 ( 
.A(n_309),
.B(n_326),
.Y(n_382)
);

AOI32xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_316),
.A3(n_319),
.B1(n_320),
.B2(n_322),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g576 ( 
.A(n_333),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_334),
.B(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_345),
.Y(n_662)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_411),
.C(n_414),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_398),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_357),
.B(n_398),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_382),
.C(n_383),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_365),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_366),
.C(n_403),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B(n_364),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_363),
.B(n_451),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_461),
.C(n_463),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_363),
.B(n_553),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_363),
.A2(n_552),
.B(n_557),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_363),
.B(n_530),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_363),
.B(n_593),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_373),
.Y(n_365)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_368),
.Y(n_531)
);

INVx3_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.C(n_396),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_385),
.B(n_434),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_388),
.A2(n_396),
.B1(n_397),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_388),
.Y(n_435)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_405),
.B(n_409),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_404),
.Y(n_399)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_402),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_404),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_412),
.C(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_406),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_415),
.A2(n_426),
.B(n_427),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_480),
.B(n_604),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_477),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_431),
.B(n_605),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_436),
.C(n_448),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_433),
.B(n_506),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_436),
.A2(n_437),
.B1(n_448),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_439),
.B(n_447),
.Y(n_437)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_447),
.B(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_465),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_465),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_454),
.B(n_460),
.Y(n_449)
);

INVx4_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_475),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_466),
.A2(n_573),
.B(n_586),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_467),
.B(n_526),
.Y(n_525)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_508),
.B(n_603),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_505),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_482),
.B(n_505),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_498),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_499),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_502),
.Y(n_664)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_563),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_532),
.B(n_562),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_511),
.B(n_513),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_528),
.C(n_529),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_514),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.Y(n_558)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_529),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_558),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_533),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_554),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_534),
.A2(n_554),
.B1(n_579),
.B2(n_580),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_534),
.Y(n_579)
);

AO221x1_ASAP7_75t_L g599 ( 
.A1(n_534),
.A2(n_554),
.B1(n_567),
.B2(n_579),
.C(n_580),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_535),
.A2(n_538),
.B(n_546),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_541),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_547),
.A2(n_550),
.B(n_552),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_554),
.Y(n_580)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_559),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_564),
.C(n_600),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_581),
.B(n_599),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_578),
.Y(n_566)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_568),
.Y(n_593)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_583),
.A2(n_589),
.B(n_598),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_585),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_584),
.B(n_585),
.Y(n_598)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_590),
.B(n_591),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_592),
.B(n_594),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_601),
.B(n_602),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_609),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_608),
.B(n_609),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_635),
.Y(n_609)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_611),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_611),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_624),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_612),
.Y(n_646)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_612),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_613),
.A2(n_615),
.B1(n_652),
.B2(n_654),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_618),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_625),
.A2(n_630),
.B1(n_631),
.B2(n_632),
.Y(n_624)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_625),
.Y(n_632)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_630),
.A2(n_631),
.B1(n_659),
.B2(n_666),
.Y(n_658)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_631),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_646),
.C(n_647),
.Y(n_645)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_635),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_639),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_641),
.B(n_674),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_R g680 ( 
.A(n_641),
.B(n_675),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_671),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_644),
.B(n_667),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_667),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_645),
.B(n_648),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_650),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_658),
.Y(n_650)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_659),
.Y(n_666)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_668),
.B(n_669),
.C(n_670),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_673),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_675),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_R g675 ( 
.A(n_676),
.B(n_678),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_677),
.Y(n_676)
);


endmodule