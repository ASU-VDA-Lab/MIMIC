module fake_jpeg_31568_n_248 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_8),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_46),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_47),
.B(n_59),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_18),
.B2(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_52),
.B1(n_57),
.B2(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_18),
.Y(n_52)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_35),
.B1(n_18),
.B2(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_31),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_27),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_35),
.A2(n_14),
.B1(n_29),
.B2(n_24),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_37),
.B1(n_40),
.B2(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_22),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_28),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_25),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_88),
.B1(n_91),
.B2(n_102),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_86),
.A2(n_100),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_42),
.B1(n_26),
.B2(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_64),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_44),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_81),
.C(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_44),
.Y(n_107)
);

INVx2_ASAP7_75t_R g109 ( 
.A(n_47),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_55),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx11_ASAP7_75t_SL g112 ( 
.A(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_60),
.B1(n_63),
.B2(n_71),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_99),
.B(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_126),
.Y(n_146)
);

XOR2x2_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_80),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_128),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_70),
.B1(n_77),
.B2(n_75),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_138),
.B1(n_99),
.B2(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_63),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_109),
.B(n_106),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_76),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_75),
.B1(n_77),
.B2(n_60),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_113),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_55),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_81),
.B1(n_61),
.B2(n_11),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_61),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_92),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_150),
.B(n_151),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_85),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_156),
.C(n_161),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_142),
.B(n_117),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_107),
.B(n_96),
.Y(n_151)
);

NAND2x1_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_94),
.C(n_90),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_90),
.B(n_92),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_164),
.B(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_131),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_127),
.C(n_12),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_95),
.B(n_113),
.C(n_11),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_130),
.B(n_12),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_82),
.B(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_108),
.Y(n_165)
);

AOI22x1_ASAP7_75t_R g166 ( 
.A1(n_139),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_118),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_157),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_135),
.B1(n_133),
.B2(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_134),
.B1(n_143),
.B2(n_123),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_123),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_152),
.B(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_184),
.B(n_167),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_130),
.B(n_129),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_129),
.C(n_10),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_162),
.C(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_190),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_159),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.C(n_194),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_155),
.B1(n_166),
.B2(n_145),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_149),
.C(n_161),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_150),
.C(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_180),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_147),
.C(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_173),
.C(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_185),
.C(n_171),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_209),
.C(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_215),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_199),
.B1(n_198),
.B2(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_222),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_194),
.B(n_190),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_182),
.B(n_213),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g228 ( 
.A(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_214),
.C(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_220),
.B1(n_224),
.B2(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_169),
.C(n_196),
.Y(n_232)
);

AO21x2_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_221),
.B(n_225),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_183),
.B(n_182),
.C(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_201),
.B1(n_182),
.B2(n_183),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_241),
.B1(n_233),
.B2(n_144),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_237),
.Y(n_245)
);

OAI221xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_233),
.B1(n_237),
.B2(n_217),
.C(n_201),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_153),
.B(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_153),
.Y(n_248)
);


endmodule