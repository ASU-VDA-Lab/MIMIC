module fake_jpeg_12877_n_85 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_30),
.B1(n_35),
.B2(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_42),
.B1(n_29),
.B2(n_26),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_27),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_33),
.C(n_12),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_60),
.C(n_10),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_67),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_11),
.B1(n_13),
.B2(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_19),
.Y(n_78)
);

OAI322xp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_69),
.A3(n_71),
.B1(n_66),
.B2(n_24),
.C1(n_20),
.C2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_76),
.C(n_74),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_77),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_73),
.Y(n_85)
);


endmodule