module fake_ariane_213_n_2126 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2126);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2126;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_2016;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_2101;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_25),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_34),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_40),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_78),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_45),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_50),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_104),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_98),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_154),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_123),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_103),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_152),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_180),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_124),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_112),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_202),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_113),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_20),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_79),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_121),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_189),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_201),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_87),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_162),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_36),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_33),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_13),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_183),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_190),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_12),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_173),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_115),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_179),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_74),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_27),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_97),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_9),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_144),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_168),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_164),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_4),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_177),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_150),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_84),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_78),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_119),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_110),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_159),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_69),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_79),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_188),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_11),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_44),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_146),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_67),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_62),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_89),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_58),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_92),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_94),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_29),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_157),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_142),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_52),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_82),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_106),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_16),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_172),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_6),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_49),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_71),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_29),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_62),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_101),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_136),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_0),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_47),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_178),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_134),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_26),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_111),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_59),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_120),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_129),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_155),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_57),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_35),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_42),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_137),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_132),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_68),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_171),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_122),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_18),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_80),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_130),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_128),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_36),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_17),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_127),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_14),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_8),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_167),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_35),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_174),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_47),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_182),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_2),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_45),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_175),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_3),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_41),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_39),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_67),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_51),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_149),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_74),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_86),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_109),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_37),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_65),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_165),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_60),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_65),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_72),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_85),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_37),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_24),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_38),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_88),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_41),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_40),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_18),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_198),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_31),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_5),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_27),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_80),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_3),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_156),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_33),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_70),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_51),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_48),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_17),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_19),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_64),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_56),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_39),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_23),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_81),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_11),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_59),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_160),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_210),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_191),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_76),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_217),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_374),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_237),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_376),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_237),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_255),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_237),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_299),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_315),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_0),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_244),
.B(n_407),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_260),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_229),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_285),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_285),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_289),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_263),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_229),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_211),
.B(n_4),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_225),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_220),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_248),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_236),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_236),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_289),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_277),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_252),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_285),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_271),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_283),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_306),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_240),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_240),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_301),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_286),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_220),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_221),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_244),
.B(n_6),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_312),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_289),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_315),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_316),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_302),
.Y(n_474)
);

BUFx2_ASAP7_75t_SL g475 ( 
.A(n_318),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_242),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_289),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_326),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_353),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_328),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_367),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_332),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_338),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_306),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_242),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_381),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_411),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_233),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_358),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_212),
.B(n_8),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_246),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_221),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_359),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_366),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_246),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_304),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_249),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_249),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_379),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_315),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_251),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_382),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_251),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_213),
.B(n_10),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_307),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_404),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_315),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_289),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_306),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_214),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_342),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_219),
.B(n_10),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_368),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_214),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_257),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_215),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_215),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_290),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_257),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_258),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_420),
.B(n_230),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_437),
.B(n_290),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_444),
.B(n_228),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_442),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_232),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_475),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_424),
.B(n_387),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_477),
.B(n_235),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_471),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_428),
.B(n_387),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_471),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_466),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_430),
.B(n_397),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_471),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_471),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_433),
.A2(n_241),
.B(n_239),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_448),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_437),
.B(n_397),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_466),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_434),
.B(n_409),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_423),
.B(n_315),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_475),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_409),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_501),
.Y(n_560)
);

BUFx8_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_429),
.B(n_438),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_501),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_512),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_501),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_423),
.B(n_346),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_512),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_468),
.B(n_253),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_511),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_436),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_440),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_455),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_422),
.B(n_231),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_511),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_438),
.B(n_253),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_511),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_518),
.Y(n_581)
);

AND3x2_ASAP7_75t_L g582 ( 
.A(n_432),
.B(n_363),
.C(n_305),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_452),
.B(n_457),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_459),
.B(n_243),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_419),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_511),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_518),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_337),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_245),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_505),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_469),
.B(n_247),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_473),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_478),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_482),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_483),
.B(n_254),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_493),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_499),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_421),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_503),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_507),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_546),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_561),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_579),
.B(n_422),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_546),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_231),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_439),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_562),
.B(n_421),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_565),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_579),
.A2(n_490),
.B1(n_516),
.B2(n_398),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_562),
.B(n_447),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_588),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_561),
.A2(n_467),
.B1(n_458),
.B2(n_461),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_592),
.B(n_425),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_588),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_531),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_592),
.B(n_425),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_569),
.A2(n_467),
.B1(n_492),
.B2(n_451),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_592),
.B(n_427),
.Y(n_632)
);

INVxp33_ASAP7_75t_SL g633 ( 
.A(n_536),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_569),
.A2(n_427),
.B1(n_472),
.B2(n_369),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_531),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_532),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_536),
.B(n_447),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_534),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_575),
.B(n_453),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_537),
.Y(n_642)
);

AND3x4_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_484),
.C(n_443),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_575),
.B(n_453),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_537),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_592),
.B(n_454),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_551),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_551),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_592),
.B(n_454),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_592),
.B(n_462),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_569),
.A2(n_380),
.B1(n_333),
.B2(n_509),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_564),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_592),
.B(n_462),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_558),
.B(n_463),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_554),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_586),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_586),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_590),
.B(n_463),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_570),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_527),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_558),
.B(n_476),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_564),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_607),
.B(n_476),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_570),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_556),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_571),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_607),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_571),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_572),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_555),
.B(n_510),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_605),
.B(n_485),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_569),
.A2(n_223),
.B1(n_224),
.B2(n_222),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_570),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_590),
.B(n_485),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_569),
.A2(n_519),
.B1(n_491),
.B2(n_497),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_573),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_573),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_605),
.B(n_491),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_570),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_590),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_570),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_561),
.A2(n_495),
.B1(n_498),
.B2(n_497),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_545),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_550),
.Y(n_688)
);

INVx11_ASAP7_75t_L g689 ( 
.A(n_561),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_545),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_590),
.B(n_495),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_561),
.B(n_498),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_590),
.B(n_502),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_550),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_550),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_588),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_590),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_598),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_587),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_526),
.B(n_502),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_553),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_550),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_587),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_588),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_526),
.B(n_504),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_588),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_528),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_606),
.B(n_504),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_574),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_556),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_553),
.B(n_513),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_526),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_555),
.B(n_305),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_574),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_582),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_555),
.A2(n_520),
.B1(n_525),
.B2(n_524),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_588),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_598),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_606),
.B(n_520),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_553),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_527),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_577),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_555),
.A2(n_598),
.B1(n_583),
.B2(n_527),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_545),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_583),
.A2(n_524),
.B1(n_525),
.B2(n_343),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_606),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_583),
.A2(n_343),
.B1(n_218),
.B2(n_266),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_587),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_528),
.B(n_426),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_606),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_583),
.B(n_343),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_606),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_527),
.A2(n_222),
.B1(n_224),
.B2(n_223),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_606),
.B(n_258),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_545),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_606),
.B(n_259),
.Y(n_742)
);

AND3x2_ASAP7_75t_L g743 ( 
.A(n_527),
.B(n_543),
.C(n_538),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_595),
.B(n_226),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_545),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_594),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_545),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_594),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_582),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_597),
.B(n_259),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_594),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_594),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_594),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_545),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_548),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_535),
.B(n_216),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_589),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_594),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_548),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_548),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_548),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_535),
.B(n_295),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_671),
.B(n_539),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_669),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_671),
.A2(n_658),
.B(n_653),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_620),
.A2(n_714),
.B1(n_725),
.B2(n_744),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_708),
.B(n_539),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_714),
.B(n_556),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_757),
.B(n_597),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_667),
.B(n_435),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_671),
.B(n_261),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_620),
.A2(n_614),
.B1(n_644),
.B2(n_641),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_671),
.B(n_261),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_763),
.B(n_599),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_649),
.B(n_599),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_650),
.B(n_603),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_723),
.B(n_262),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_618),
.B(n_604),
.C(n_603),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_733),
.B(n_604),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_714),
.B(n_556),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_627),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_669),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_676),
.B(n_608),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_691),
.B(n_608),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_723),
.B(n_262),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_633),
.B(n_445),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_693),
.B(n_610),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_635),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_723),
.B(n_362),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_758),
.B(n_744),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_723),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_625),
.B(n_362),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_758),
.B(n_610),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_630),
.B(n_399),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_678),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_621),
.B(n_456),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_613),
.B(n_595),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_612),
.B(n_464),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_674),
.A2(n_591),
.B1(n_596),
.B2(n_585),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_663),
.B(n_474),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_702),
.B(n_595),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_635),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_637),
.B(n_479),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_683),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_661),
.B(n_481),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_714),
.A2(n_600),
.B1(n_609),
.B2(n_602),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_721),
.B(n_600),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_611),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_632),
.B(n_600),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_713),
.B(n_602),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_713),
.B(n_602),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_646),
.B(n_399),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_654),
.B(n_227),
.C(n_226),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_722),
.B(n_609),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_701),
.B(n_609),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_623),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_619),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_636),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_672),
.B(n_486),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_683),
.B(n_415),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_714),
.A2(n_589),
.B1(n_594),
.B2(n_593),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_680),
.B(n_487),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_619),
.Y(n_830)
);

AND2x6_ASAP7_75t_L g831 ( 
.A(n_688),
.B(n_308),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_674),
.A2(n_591),
.B1(n_596),
.B2(n_585),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_714),
.A2(n_589),
.B1(n_593),
.B2(n_581),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_706),
.B(n_601),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_686),
.Y(n_835)
);

NAND2x1_ASAP7_75t_L g836 ( 
.A(n_665),
.B(n_549),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_683),
.B(n_415),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_670),
.B(n_601),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_686),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_617),
.B(n_488),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_612),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_615),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_615),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_655),
.B(n_538),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_670),
.B(n_578),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_743),
.B(n_538),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_636),
.Y(n_847)
);

BUFx6f_ASAP7_75t_SL g848 ( 
.A(n_750),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_670),
.B(n_578),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_688),
.A2(n_581),
.B(n_567),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_670),
.B(n_543),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_636),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_750),
.B(n_543),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_547),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_622),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_496),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_SL g857 ( 
.A(n_613),
.B(n_227),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_655),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_699),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_662),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_662),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_716),
.B(n_547),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_662),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_735),
.B(n_547),
.Y(n_864)
);

AND2x6_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_308),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_638),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_622),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_714),
.B(n_593),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_659),
.A2(n_587),
.B(n_533),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_712),
.B(n_506),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_731),
.A2(n_559),
.B1(n_360),
.B2(n_347),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_642),
.B(n_559),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_683),
.B(n_416),
.Y(n_873)
);

NOR2x1p5_ASAP7_75t_L g874 ( 
.A(n_656),
.B(n_234),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_638),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_712),
.B(n_515),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_698),
.B(n_416),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_642),
.B(n_559),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_698),
.B(n_623),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_645),
.B(n_393),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_639),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_682),
.Y(n_882)
);

AND3x1_ASAP7_75t_L g883 ( 
.A(n_728),
.B(n_238),
.C(n_234),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_645),
.B(n_417),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_651),
.A2(n_360),
.B1(n_371),
.B2(n_331),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_639),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_629),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_648),
.A2(n_293),
.B(n_375),
.C(n_377),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_682),
.B(n_517),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_659),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_698),
.B(n_417),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_629),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_648),
.B(n_264),
.Y(n_893)
);

AO22x2_ASAP7_75t_L g894 ( 
.A1(n_643),
.A2(n_371),
.B1(n_354),
.B2(n_331),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_657),
.A2(n_355),
.B1(n_238),
.B2(n_250),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_698),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_623),
.B(n_256),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_652),
.B(n_265),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_652),
.B(n_272),
.Y(n_899)
);

OAI22xp33_ASAP7_75t_L g900 ( 
.A1(n_738),
.A2(n_383),
.B1(n_250),
.B2(n_351),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_623),
.B(n_270),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_640),
.B(n_273),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_640),
.B(n_647),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_647),
.B(n_274),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_716),
.B(n_351),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_717),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_710),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_666),
.B(n_275),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_715),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_660),
.B(n_352),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_666),
.B(n_276),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_660),
.B(n_356),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_692),
.A2(n_300),
.B1(n_298),
.B2(n_364),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_660),
.B(n_361),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_623),
.B(n_556),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_751),
.B(n_365),
.C(n_361),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_715),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_738),
.B(n_365),
.Y(n_919)
);

AO221x1_ASAP7_75t_L g920 ( 
.A1(n_643),
.A2(n_346),
.B1(n_385),
.B2(n_389),
.C(n_278),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_685),
.B(n_288),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_699),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_623),
.B(n_296),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_666),
.B(n_279),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_660),
.B(n_370),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_724),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_677),
.B(n_370),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_626),
.B(n_311),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_724),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_634),
.B(n_373),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_727),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_668),
.B(n_282),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_626),
.B(n_314),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_668),
.B(n_294),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_631),
.B(n_383),
.C(n_373),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_814),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_842),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_775),
.B(n_643),
.Y(n_938)
);

AOI21xp33_ASAP7_75t_L g939 ( 
.A1(n_930),
.A2(n_624),
.B(n_699),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_804),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_766),
.A2(n_664),
.B(n_659),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_764),
.A2(n_673),
.B(n_668),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_768),
.A2(n_679),
.B(n_673),
.C(n_727),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_834),
.B(n_719),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_SL g945 ( 
.A1(n_774),
.A2(n_679),
.B(n_673),
.C(n_730),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_838),
.B(n_719),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_773),
.B(n_679),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_844),
.B(n_841),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_786),
.A2(n_792),
.B(n_787),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_821),
.B(n_719),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_843),
.B(n_700),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_771),
.B(n_659),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_858),
.B(n_384),
.Y(n_953)
);

O2A1O1Ixp5_ASAP7_75t_L g954 ( 
.A1(n_797),
.A2(n_742),
.B(n_740),
.C(n_734),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_919),
.A2(n_906),
.B(n_900),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_823),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_664),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_822),
.A2(n_703),
.B(n_694),
.C(n_695),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_764),
.A2(n_734),
.B(n_730),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_850),
.A2(n_737),
.B(n_729),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_805),
.B(n_832),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_889),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_862),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_778),
.A2(n_675),
.B(n_664),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_779),
.A2(n_675),
.B(n_664),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_889),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_882),
.B(n_700),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_782),
.B(n_675),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_862),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_815),
.A2(n_681),
.B(n_675),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_769),
.B(n_681),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_774),
.A2(n_684),
.B(n_681),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_862),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_784),
.A2(n_737),
.B(n_729),
.Y(n_974)
);

CKINVDCx6p67_ASAP7_75t_R g975 ( 
.A(n_848),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_776),
.A2(n_684),
.B(n_681),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_846),
.B(n_665),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_907),
.B(n_386),
.C(n_384),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_848),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_795),
.B(n_684),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_776),
.A2(n_684),
.B(n_709),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_789),
.A2(n_696),
.B(n_695),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_854),
.A2(n_720),
.B(n_700),
.C(n_704),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_823),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_864),
.B(n_696),
.Y(n_985)
);

CKINVDCx10_ASAP7_75t_R g986 ( 
.A(n_848),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_824),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_879),
.A2(n_703),
.B(n_705),
.Y(n_988)
);

OAI321xp33_ASAP7_75t_L g989 ( 
.A1(n_927),
.A2(n_317),
.A3(n_330),
.B1(n_335),
.B2(n_378),
.C(n_357),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_796),
.B(n_626),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_796),
.B(n_626),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_807),
.B(n_700),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_895),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_879),
.A2(n_707),
.B(n_705),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_827),
.A2(n_873),
.B(n_877),
.C(n_837),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_883),
.A2(n_616),
.B1(n_759),
.B2(n_754),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_904),
.A2(n_718),
.B(n_707),
.Y(n_997)
);

NOR2x1_ASAP7_75t_R g998 ( 
.A(n_772),
.B(n_927),
.Y(n_998)
);

AOI33xp33_ASAP7_75t_L g999 ( 
.A1(n_765),
.A2(n_396),
.A3(n_418),
.B1(n_414),
.B2(n_412),
.B3(n_410),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_827),
.A2(n_718),
.B(n_747),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_813),
.B(n_704),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_830),
.A2(n_704),
.B(n_732),
.C(n_739),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_846),
.B(n_689),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_853),
.B(n_704),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_853),
.B(n_732),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_855),
.A2(n_739),
.B1(n_732),
.B2(n_736),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_837),
.A2(n_749),
.B(n_747),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_772),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_867),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_873),
.A2(n_891),
.B(n_877),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_791),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_840),
.B(n_388),
.C(n_386),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_853),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_790),
.B(n_665),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_887),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_891),
.A2(n_799),
.B(n_797),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_894),
.A2(n_616),
.B1(n_759),
.B2(n_754),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_870),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_890),
.B(n_626),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_894),
.A2(n_616),
.B1(n_665),
.B2(n_711),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_856),
.B(n_388),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_892),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_785),
.A2(n_732),
.B(n_739),
.C(n_749),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_890),
.B(n_626),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_851),
.B(n_739),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_799),
.A2(n_753),
.B(n_752),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_823),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_791),
.A2(n_808),
.B(n_793),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_818),
.A2(n_753),
.B(n_752),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_845),
.B(n_616),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_818),
.A2(n_736),
.B(n_690),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_849),
.B(n_616),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_823),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_793),
.A2(n_736),
.B(n_690),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_800),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_874),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_808),
.A2(n_690),
.B(n_687),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_825),
.A2(n_726),
.B(n_687),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_890),
.B(n_697),
.Y(n_1039)
);

OAI21xp33_ASAP7_75t_SL g1040 ( 
.A1(n_801),
.A2(n_711),
.B(n_687),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_901),
.A2(n_410),
.B(n_392),
.C(n_394),
.Y(n_1041)
);

AO21x1_ASAP7_75t_L g1042 ( 
.A1(n_780),
.A2(n_794),
.B(n_788),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_825),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_802),
.B(n_394),
.C(n_392),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_880),
.B(n_616),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_847),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_846),
.B(n_697),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_767),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_767),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_835),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_810),
.B(n_697),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_847),
.A2(n_741),
.B(n_726),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_868),
.A2(n_741),
.B(n_726),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_908),
.A2(n_697),
.B1(n_395),
.B2(n_396),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_852),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_910),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_798),
.B(n_616),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_876),
.B(n_395),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_918),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_820),
.B(n_697),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_897),
.A2(n_923),
.B(n_902),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_810),
.B(n_697),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_772),
.B(n_711),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_806),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_780),
.A2(n_354),
.B(n_741),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_894),
.A2(n_711),
.B1(n_327),
.B2(n_303),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_835),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_781),
.B(n_400),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_911),
.B(n_400),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_926),
.A2(n_931),
.B1(n_929),
.B2(n_872),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_852),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_935),
.B(n_913),
.Y(n_1072)
);

CKINVDCx10_ASAP7_75t_R g1073 ( 
.A(n_826),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_829),
.B(n_401),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_915),
.B(n_925),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_770),
.B(n_346),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_788),
.A2(n_762),
.B(n_761),
.C(n_760),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_809),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_860),
.A2(n_746),
.B(n_745),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_860),
.A2(n_746),
.B(n_745),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_878),
.A2(n_408),
.B1(n_401),
.B2(n_403),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_861),
.A2(n_746),
.B(n_745),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_839),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_861),
.A2(n_755),
.B(n_748),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_869),
.A2(n_755),
.B(n_748),
.Y(n_1085)
);

OAI321xp33_ASAP7_75t_L g1086 ( 
.A1(n_871),
.A2(n_389),
.A3(n_346),
.B1(n_385),
.B2(n_533),
.C(n_541),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_863),
.A2(n_755),
.B(n_748),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_816),
.B(n_403),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_896),
.B(n_839),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_863),
.A2(n_896),
.B(n_794),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_888),
.A2(n_406),
.B(n_414),
.C(n_412),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_866),
.A2(n_762),
.B(n_761),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_859),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_866),
.A2(n_762),
.B(n_761),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_817),
.B(n_406),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_875),
.A2(n_886),
.B(n_881),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_819),
.B(n_418),
.C(n_408),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_875),
.A2(n_756),
.B(n_760),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_811),
.B(n_756),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_859),
.B(n_756),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_893),
.B(n_760),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_898),
.B(n_309),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_922),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_899),
.B(n_310),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_884),
.B(n_319),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_833),
.B(n_903),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_886),
.A2(n_628),
.B(n_529),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_885),
.A2(n_324),
.B(n_325),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_917),
.B(n_329),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_905),
.B(n_336),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_909),
.B(n_345),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_912),
.A2(n_529),
.B(n_533),
.C(n_541),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_924),
.B(n_13),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_L g1114 ( 
.A(n_803),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_L g1115 ( 
.A(n_831),
.B(n_628),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_932),
.B(n_14),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_836),
.A2(n_628),
.B(n_529),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_934),
.A2(n_628),
.B(n_541),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_922),
.A2(n_628),
.B(n_542),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_770),
.A2(n_628),
.B(n_542),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_914),
.B(n_15),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_783),
.A2(n_542),
.B(n_580),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_921),
.B(n_267),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_783),
.A2(n_552),
.B(n_580),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_936),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_938),
.A2(n_812),
.B(n_857),
.C(n_923),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_961),
.B(n_831),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1085),
.A2(n_933),
.B(n_928),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_938),
.A2(n_933),
.B(n_928),
.C(n_902),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_952),
.B(n_831),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1048),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_962),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1048),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_937),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1048),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_949),
.A2(n_803),
.B(n_916),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_971),
.A2(n_803),
.B(n_916),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_987),
.Y(n_1138)
);

AO32x1_ASAP7_75t_L g1139 ( 
.A1(n_1070),
.A2(n_552),
.A3(n_563),
.B1(n_566),
.B2(n_576),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1075),
.A2(n_897),
.B(n_920),
.C(n_865),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_940),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_952),
.B(n_831),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_957),
.B(n_831),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1002),
.A2(n_865),
.B(n_831),
.C(n_576),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_955),
.A2(n_828),
.B1(n_339),
.B2(n_334),
.C(n_269),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_937),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_971),
.A2(n_803),
.B(n_865),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1069),
.A2(n_552),
.B(n_563),
.C(n_566),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1048),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_940),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_973),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_977),
.B(n_865),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1072),
.B(n_268),
.C(n_280),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1018),
.A2(n_865),
.B1(n_281),
.B2(n_350),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1076),
.A2(n_865),
.B1(n_323),
.B2(n_321),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_969),
.B(n_284),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_SL g1158 ( 
.A1(n_993),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1104),
.A2(n_563),
.B(n_566),
.C(n_576),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_969),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_956),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1064),
.B(n_297),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1068),
.A2(n_313),
.B(n_320),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_977),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1008),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1009),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_986),
.B(n_340),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1011),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1014),
.B(n_341),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1078),
.B(n_963),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_947),
.B(n_948),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1114),
.B(n_344),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_963),
.B(n_580),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_950),
.A2(n_349),
.B(n_346),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1103),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_950),
.A2(n_385),
.B(n_389),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_957),
.B(n_556),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1114),
.B(n_530),
.Y(n_1178)
);

OAI21xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1076),
.A2(n_15),
.B(n_16),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1008),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1050),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_956),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1074),
.B(n_19),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1015),
.Y(n_1184)
);

BUFx4f_ASAP7_75t_L g1185 ( 
.A(n_975),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1072),
.B(n_530),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_944),
.A2(n_385),
.B(n_389),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1104),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_964),
.A2(n_385),
.B(n_389),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_965),
.A2(n_584),
.B(n_548),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_SL g1192 ( 
.A(n_998),
.B(n_556),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1091),
.A2(n_22),
.B(n_26),
.C(n_28),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_1058),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_1003),
.B(n_549),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_985),
.B(n_556),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_956),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1022),
.B(n_556),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1091),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1010),
.A2(n_549),
.B(n_530),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_941),
.A2(n_584),
.B(n_548),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1021),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1063),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1035),
.B(n_567),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_978),
.A2(n_32),
.B(n_34),
.C(n_38),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1056),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1036),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1059),
.A2(n_549),
.B1(n_42),
.B2(n_43),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_968),
.A2(n_584),
.B(n_548),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_970),
.A2(n_584),
.B(n_548),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1012),
.B(n_557),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1113),
.A2(n_584),
.B(n_560),
.C(n_557),
.Y(n_1212)
);

BUFx8_ASAP7_75t_L g1213 ( 
.A(n_953),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_995),
.A2(n_584),
.B(n_560),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1043),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_979),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1013),
.B(n_1106),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1113),
.A2(n_584),
.B(n_560),
.C(n_557),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1053),
.A2(n_567),
.B(n_549),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_939),
.B(n_32),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1102),
.A2(n_1105),
.B(n_1116),
.C(n_1121),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1073),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1046),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1116),
.A2(n_549),
.B1(n_44),
.B2(n_46),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_951),
.B(n_43),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1055),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1013),
.B(n_567),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1121),
.A2(n_584),
.B(n_560),
.C(n_557),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_L g1229 ( 
.A(n_956),
.B(n_567),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1109),
.A2(n_567),
.B1(n_48),
.B2(n_49),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1071),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1095),
.B(n_46),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_967),
.B(n_50),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_L g1234 ( 
.A(n_984),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_946),
.B(n_567),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1050),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1004),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_995),
.A2(n_560),
.B(n_557),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1067),
.Y(n_1239)
);

BUFx8_ASAP7_75t_SL g1240 ( 
.A(n_984),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1044),
.B(n_530),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_980),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1005),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1067),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1063),
.B(n_530),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_L g1246 ( 
.A(n_1097),
.B(n_53),
.C(n_54),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1101),
.A2(n_560),
.B(n_557),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1110),
.B(n_56),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1049),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1083),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1016),
.A2(n_560),
.B(n_540),
.C(n_544),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1047),
.B(n_1025),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_984),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_943),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_1254)
);

CKINVDCx14_ASAP7_75t_R g1255 ( 
.A(n_1003),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1049),
.Y(n_1256)
);

OR2x6_ASAP7_75t_SL g1257 ( 
.A(n_1081),
.B(n_61),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1090),
.A2(n_567),
.B(n_126),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1095),
.B(n_63),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_984),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_981),
.A2(n_560),
.B(n_557),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_943),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1111),
.A2(n_66),
.B(n_72),
.C(n_73),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_544),
.B(n_540),
.C(n_530),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1047),
.B(n_544),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1088),
.B(n_73),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1093),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1108),
.B(n_75),
.Y(n_1268)
);

BUFx4f_ASAP7_75t_L g1269 ( 
.A(n_1027),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1066),
.A2(n_544),
.B(n_540),
.C(n_530),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1093),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1083),
.B(n_544),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1027),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1020),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_958),
.B(n_992),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_958),
.B(n_567),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1099),
.B(n_567),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1027),
.Y(n_1278)
);

NAND3xp33_ASAP7_75t_SL g1279 ( 
.A(n_999),
.B(n_77),
.C(n_83),
.Y(n_1279)
);

OAI21xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1019),
.A2(n_91),
.B(n_95),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1100),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1096),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1001),
.B(n_544),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1027),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1033),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_994),
.A2(n_960),
.B(n_945),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1220),
.A2(n_1020),
.B1(n_1042),
.B2(n_1123),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1251),
.A2(n_1065),
.A3(n_1002),
.B(n_1031),
.Y(n_1288)
);

BUFx4f_ASAP7_75t_L g1289 ( 
.A(n_1132),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1136),
.A2(n_1115),
.B(n_945),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1257),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1130),
.A2(n_1040),
.B(n_1024),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1160),
.B(n_1033),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1125),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1130),
.A2(n_1019),
.B(n_1024),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1160),
.B(n_1164),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1221),
.A2(n_1057),
.B(n_942),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1142),
.A2(n_1039),
.B(n_974),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_988),
.B(n_997),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1164),
.B(n_1150),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1248),
.A2(n_1086),
.B(n_1045),
.C(n_1017),
.Y(n_1301)
);

CKINVDCx12_ASAP7_75t_R g1302 ( 
.A(n_1230),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1266),
.A2(n_954),
.B(n_1041),
.C(n_983),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1156),
.B(n_1030),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1183),
.A2(n_1041),
.B(n_1023),
.C(n_1054),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1171),
.B(n_982),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1134),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1194),
.B(n_1089),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1146),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1222),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1141),
.B(n_1033),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1166),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1147),
.A2(n_1028),
.B(n_1000),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1184),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1234),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1213),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1142),
.A2(n_1032),
.B(n_972),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1219),
.A2(n_1092),
.B(n_1094),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1170),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1143),
.A2(n_1039),
.B(n_1051),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1167),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1268),
.A2(n_996),
.B(n_1077),
.C(n_1026),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1206),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1188),
.B(n_1029),
.C(n_1112),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1252),
.B(n_1060),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1286),
.A2(n_1201),
.B(n_1128),
.Y(n_1327)
);

OAI21xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1232),
.A2(n_990),
.B(n_991),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1238),
.A2(n_1098),
.B(n_1052),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1143),
.A2(n_1051),
.B(n_1062),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1137),
.A2(n_1062),
.B(n_990),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1191),
.B(n_1089),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1202),
.B(n_1033),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1275),
.A2(n_991),
.B(n_976),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1275),
.A2(n_1006),
.B(n_1034),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1252),
.A2(n_1007),
.B(n_959),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1151),
.B(n_1080),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1156),
.A2(n_1100),
.B(n_1087),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1144),
.A2(n_1084),
.B(n_1037),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1259),
.A2(n_1118),
.B(n_1038),
.C(n_1079),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1127),
.A2(n_1082),
.B(n_1122),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1255),
.A2(n_1120),
.B1(n_1119),
.B2(n_1124),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1181),
.B(n_1061),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1129),
.A2(n_1107),
.B(n_1117),
.C(n_544),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1127),
.A2(n_540),
.B(n_100),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1247),
.A2(n_540),
.B(n_105),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1191),
.B(n_99),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1126),
.A2(n_540),
.B(n_114),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1217),
.B(n_540),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1228),
.A2(n_107),
.B(n_116),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1214),
.A2(n_117),
.B(n_118),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1196),
.A2(n_125),
.B(n_133),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1274),
.A2(n_138),
.B1(n_143),
.B2(n_147),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1211),
.A2(n_153),
.B(n_170),
.C(n_187),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1203),
.B(n_192),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1181),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1212),
.A2(n_193),
.B(n_194),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1261),
.A2(n_1190),
.B(n_1210),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1155),
.B(n_195),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1177),
.A2(n_197),
.B(n_204),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1177),
.A2(n_1218),
.B(n_1283),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1179),
.A2(n_207),
.B(n_1205),
.C(n_1163),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1270),
.A2(n_1258),
.A3(n_1282),
.B(n_1187),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_SL g1364 ( 
.A1(n_1224),
.A2(n_1241),
.B(n_1254),
.C(n_1262),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_L g1365 ( 
.A(n_1250),
.B(n_1236),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1283),
.A2(n_1189),
.B(n_1209),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1176),
.A2(n_1186),
.B(n_1276),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1224),
.A2(n_1254),
.B(n_1262),
.C(n_1157),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1168),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1217),
.B(n_1237),
.Y(n_1370)
);

AO32x2_ASAP7_75t_L g1371 ( 
.A1(n_1242),
.A2(n_1208),
.A3(n_1139),
.B1(n_1199),
.B2(n_1193),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1196),
.A2(n_1235),
.B(n_1152),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1235),
.A2(n_1152),
.B(n_1245),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1213),
.B(n_1239),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1243),
.B(n_1203),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1276),
.A2(n_1204),
.B(n_1198),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1152),
.A2(n_1269),
.B(n_1234),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1240),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1263),
.A2(n_1225),
.B(n_1233),
.C(n_1153),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1215),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1198),
.A2(n_1204),
.B(n_1159),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1264),
.A2(n_1140),
.B(n_1174),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1246),
.B(n_1242),
.C(n_1145),
.Y(n_1383)
);

OAI22x1_ASAP7_75t_L g1384 ( 
.A1(n_1244),
.A2(n_1172),
.B1(n_1162),
.B2(n_1154),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1148),
.A2(n_1281),
.B(n_1265),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1280),
.A2(n_1208),
.B(n_1169),
.C(n_1279),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1269),
.A2(n_1272),
.B(n_1139),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1132),
.Y(n_1388)
);

NOR4xp25_ASAP7_75t_L g1389 ( 
.A(n_1249),
.B(n_1256),
.C(n_1267),
.D(n_1178),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1271),
.A2(n_1216),
.B(n_1250),
.C(n_1175),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1207),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1158),
.B(n_1207),
.Y(n_1392)
);

AOI221x1_ASAP7_75t_L g1393 ( 
.A1(n_1227),
.A2(n_1223),
.B1(n_1226),
.B2(n_1231),
.C(n_1173),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1139),
.A2(n_1284),
.B(n_1277),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1131),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1173),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1277),
.A2(n_1229),
.B(n_1180),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1165),
.A2(n_1161),
.B(n_1278),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1285),
.B(n_1131),
.Y(n_1399)
);

BUFx8_ASAP7_75t_L g1400 ( 
.A(n_1131),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1133),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1161),
.A2(n_1278),
.B(n_1273),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1133),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1161),
.A2(n_1278),
.B(n_1273),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1192),
.A2(n_1185),
.B(n_1135),
.C(n_1149),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1182),
.B(n_1273),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1182),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1197),
.B(n_1253),
.Y(n_1409)
);

NOR2x1_ASAP7_75t_SL g1410 ( 
.A(n_1195),
.B(n_1197),
.Y(n_1410)
);

BUFx8_ASAP7_75t_L g1411 ( 
.A(n_1197),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1253),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1253),
.A2(n_1260),
.B(n_1195),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1260),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1260),
.A2(n_1195),
.B(n_1192),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1185),
.A2(n_775),
.B(n_1221),
.C(n_961),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1221),
.A2(n_938),
.B(n_775),
.C(n_1248),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1251),
.A2(n_1065),
.A3(n_1042),
.B(n_1270),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1221),
.A2(n_961),
.B(n_775),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1194),
.B(n_948),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1125),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1160),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1221),
.A2(n_938),
.B(n_775),
.C(n_1248),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1252),
.B(n_961),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1221),
.B(n_775),
.C(n_961),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1125),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1132),
.Y(n_1432)
);

BUFx12f_ASAP7_75t_L g1433 ( 
.A(n_1222),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1252),
.B(n_961),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1125),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1222),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1441)
);

OR2x6_ASAP7_75t_L g1442 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1200),
.A2(n_1219),
.B(n_1286),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1183),
.A2(n_961),
.B1(n_938),
.B2(n_775),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1171),
.B(n_667),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1240),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1125),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1125),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1194),
.B(n_657),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1252),
.B(n_961),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1251),
.A2(n_1065),
.A3(n_1042),
.B(n_1270),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1220),
.A2(n_938),
.B1(n_876),
.B2(n_870),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1134),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1136),
.A2(n_949),
.B(n_961),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1343),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1454),
.A2(n_1446),
.B1(n_1383),
.B2(n_1430),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1289),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1446),
.A2(n_1353),
.B1(n_1348),
.B2(n_1302),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1353),
.A2(n_1417),
.B1(n_1427),
.B2(n_1392),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1423),
.B(n_1320),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1400),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1422),
.A2(n_1291),
.B1(n_1348),
.B2(n_1287),
.Y(n_1464)
);

BUFx8_ASAP7_75t_SL g1465 ( 
.A(n_1311),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1294),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_1434),
.B2(n_1428),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1305),
.A2(n_1350),
.B1(n_1328),
.B2(n_1347),
.Y(n_1468)
);

BUFx2_ASAP7_75t_SL g1469 ( 
.A(n_1378),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1379),
.A2(n_1416),
.B1(n_1428),
.B2(n_1452),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1434),
.A2(n_1386),
.B1(n_1362),
.B2(n_1308),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1411),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1305),
.A2(n_1350),
.B1(n_1359),
.B2(n_1368),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1420),
.A2(n_1436),
.B(n_1425),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1309),
.A2(n_1370),
.B1(n_1451),
.B2(n_1382),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1384),
.A2(n_1370),
.B1(n_1447),
.B2(n_1356),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1411),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1304),
.A2(n_1310),
.B1(n_1455),
.B2(n_1306),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1289),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1433),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1378),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1382),
.A2(n_1352),
.B1(n_1374),
.B2(n_1364),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1440),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1303),
.Y(n_1484)
);

BUFx4f_ASAP7_75t_L g1485 ( 
.A(n_1378),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1307),
.A2(n_1375),
.B1(n_1439),
.B2(n_1442),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1337),
.A2(n_1313),
.B1(n_1450),
.B2(n_1449),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1448),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1332),
.A2(n_1442),
.B1(n_1296),
.B2(n_1365),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1315),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1400),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1324),
.A2(n_1424),
.B1(n_1431),
.B2(n_1437),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1369),
.A2(n_1380),
.B1(n_1326),
.B2(n_1375),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1399),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1333),
.A2(n_1301),
.B1(n_1426),
.B2(n_1323),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1401),
.Y(n_1496)
);

BUFx12f_ASAP7_75t_L g1497 ( 
.A(n_1448),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1448),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1326),
.A2(n_1396),
.B1(n_1442),
.B2(n_1317),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1296),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1322),
.Y(n_1501)
);

BUFx12f_ASAP7_75t_L g1502 ( 
.A(n_1391),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1388),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1432),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1300),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1297),
.A2(n_1376),
.B1(n_1300),
.B2(n_1325),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1352),
.A2(n_1357),
.B1(n_1410),
.B2(n_1297),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1403),
.B(n_1408),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1412),
.Y(n_1509)
);

CKINVDCx11_ASAP7_75t_R g1510 ( 
.A(n_1406),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1414),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1357),
.A2(n_1371),
.B1(n_1397),
.B2(n_1312),
.Y(n_1512)
);

CKINVDCx11_ASAP7_75t_R g1513 ( 
.A(n_1406),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1376),
.A2(n_1318),
.B1(n_1456),
.B2(n_1441),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1371),
.A2(n_1312),
.B1(n_1377),
.B2(n_1415),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1390),
.A2(n_1438),
.B1(n_1443),
.B2(n_1316),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1407),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1371),
.A2(n_1373),
.B1(n_1290),
.B2(n_1345),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1318),
.A2(n_1372),
.B1(n_1381),
.B2(n_1298),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1314),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1293),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1406),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1349),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1381),
.A2(n_1349),
.B1(n_1355),
.B2(n_1336),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1413),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1342),
.A2(n_1316),
.B1(n_1330),
.B2(n_1335),
.Y(n_1526)
);

INVx3_ASAP7_75t_SL g1527 ( 
.A(n_1395),
.Y(n_1527)
);

INVx6_ASAP7_75t_L g1528 ( 
.A(n_1405),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_L g1529 ( 
.A(n_1367),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1331),
.A2(n_1321),
.B1(n_1292),
.B2(n_1338),
.Y(n_1530)
);

CKINVDCx16_ASAP7_75t_R g1531 ( 
.A(n_1389),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1367),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1402),
.Y(n_1533)
);

INVx6_ASAP7_75t_L g1534 ( 
.A(n_1409),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1295),
.A2(n_1314),
.B1(n_1334),
.B2(n_1394),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1360),
.A2(n_1361),
.B1(n_1341),
.B2(n_1387),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1393),
.A2(n_1398),
.B1(n_1404),
.B2(n_1339),
.Y(n_1537)
);

INVx3_ASAP7_75t_SL g1538 ( 
.A(n_1389),
.Y(n_1538)
);

INVx6_ASAP7_75t_L g1539 ( 
.A(n_1354),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1385),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1340),
.A2(n_1344),
.B1(n_1366),
.B2(n_1346),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1363),
.A2(n_1453),
.B1(n_1419),
.B2(n_1351),
.Y(n_1542)
);

INVx8_ASAP7_75t_L g1543 ( 
.A(n_1419),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1319),
.B(n_1299),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1329),
.A2(n_1421),
.B1(n_1444),
.B2(n_1435),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1327),
.A2(n_1418),
.B1(n_1429),
.B2(n_1445),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1363),
.A2(n_1453),
.B1(n_1288),
.B2(n_1358),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1363),
.B(n_1453),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1288),
.A2(n_938),
.B1(n_1446),
.B2(n_1427),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1294),
.Y(n_1550)
);

BUFx12f_ASAP7_75t_L g1551 ( 
.A(n_1311),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1433),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1289),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1294),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1555)
);

OAI22x1_ASAP7_75t_SL g1556 ( 
.A1(n_1311),
.A2(n_657),
.B1(n_656),
.B2(n_1222),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_894),
.B2(n_426),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_894),
.B2(n_426),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1446),
.A2(n_961),
.B1(n_938),
.B2(n_620),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1343),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1294),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1311),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1400),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1294),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1566)
);

OR2x6_ASAP7_75t_L g1567 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1311),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1400),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1423),
.B(n_1320),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1343),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1573)
);

CKINVDCx6p67_ASAP7_75t_R g1574 ( 
.A(n_1433),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1423),
.B(n_1320),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1411),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1423),
.B(n_1320),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_894),
.B2(n_426),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1400),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1581)
);

CKINVDCx11_ASAP7_75t_R g1582 ( 
.A(n_1433),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1433),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1294),
.Y(n_1585)
);

OAI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1446),
.A2(n_961),
.B1(n_938),
.B2(n_620),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1400),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1400),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_894),
.B2(n_426),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1433),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_1433),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1596)
);

CKINVDCx6p67_ASAP7_75t_R g1597 ( 
.A(n_1433),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1423),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_1427),
.B2(n_1417),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1311),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1294),
.Y(n_1604)
);

INVx5_ASAP7_75t_L g1605 ( 
.A(n_1439),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1417),
.A2(n_1427),
.B(n_938),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_1427),
.B2(n_1417),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1294),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1294),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_1427),
.B2(n_1417),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1454),
.A2(n_938),
.B1(n_1446),
.B2(n_894),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1343),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1446),
.A2(n_938),
.B1(n_1427),
.B2(n_1417),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1311),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1400),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1457),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1457),
.B(n_1561),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1561),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1460),
.A2(n_1464),
.B1(n_1579),
.B2(n_1558),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1571),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1473),
.A2(n_1530),
.B(n_1474),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1525),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1529),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1464),
.A2(n_1590),
.B1(n_1557),
.B2(n_1559),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1466),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1520),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1523),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1531),
.B(n_1487),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1541),
.A2(n_1544),
.B(n_1536),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1525),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1504),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1529),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1484),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1520),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1490),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1487),
.B(n_1549),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1550),
.B(n_1554),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1559),
.A2(n_1586),
.B1(n_1589),
.B2(n_1555),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1544),
.A2(n_1536),
.B(n_1546),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1525),
.B(n_1533),
.Y(n_1642)
);

NAND2x1_ASAP7_75t_L g1643 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1546),
.A2(n_1535),
.B(n_1514),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1538),
.B(n_1548),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1562),
.B(n_1565),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1585),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1604),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1492),
.B(n_1519),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1532),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1532),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1461),
.A2(n_1607),
.B(n_1600),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1492),
.B(n_1467),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1586),
.A2(n_1612),
.B1(n_1615),
.B2(n_1470),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1535),
.A2(n_1514),
.B(n_1545),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1556),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1467),
.B(n_1576),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1583),
.B(n_1596),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1540),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1522),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1603),
.B(n_1494),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1543),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1471),
.A2(n_1495),
.A3(n_1478),
.B(n_1496),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1525),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1482),
.B(n_1468),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1524),
.A2(n_1506),
.B(n_1499),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1465),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1458),
.B(n_1606),
.C(n_1475),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1539),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1508),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1458),
.A2(n_1591),
.B1(n_1581),
.B2(n_1592),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1462),
.B(n_1570),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1547),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1509),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1575),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1493),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1517),
.B(n_1599),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1539),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1493),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1472),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1511),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1528),
.A2(n_1581),
.B1(n_1613),
.B2(n_1609),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1526),
.Y(n_1685)
);

OAI22x1_ASAP7_75t_L g1686 ( 
.A1(n_1538),
.A2(n_1489),
.B1(n_1476),
.B2(n_1605),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1526),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1528),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1486),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1528),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1578),
.B(n_1506),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1486),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1542),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1542),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1567),
.A2(n_1595),
.B1(n_1613),
.B2(n_1609),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1537),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1539),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1537),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1512),
.A2(n_1518),
.B(n_1507),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1534),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1472),
.Y(n_1701)
);

INVxp33_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1515),
.B(n_1524),
.Y(n_1703)
);

BUFx12f_ASAP7_75t_L g1704 ( 
.A(n_1498),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1555),
.B(n_1560),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1476),
.B(n_1499),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1616),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1521),
.A2(n_1608),
.B(n_1566),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1527),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1560),
.A2(n_1608),
.B(n_1573),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1566),
.A2(n_1589),
.B1(n_1573),
.B2(n_1602),
.Y(n_1711)
);

AO21x1_ASAP7_75t_L g1712 ( 
.A1(n_1572),
.A2(n_1602),
.B(n_1595),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1572),
.B(n_1598),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1591),
.B(n_1598),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1534),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1500),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1527),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1592),
.B(n_1505),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1513),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1472),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1477),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1463),
.A2(n_1580),
.B(n_1503),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1459),
.B(n_1617),
.Y(n_1723)
);

NAND2x1p5_ASAP7_75t_L g1724 ( 
.A(n_1479),
.B(n_1553),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1477),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1502),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1491),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1491),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1491),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1577),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1577),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1564),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1621),
.A2(n_1626),
.B1(n_1670),
.B2(n_1640),
.C(n_1667),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1691),
.B(n_1651),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1691),
.B(n_1651),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1635),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1670),
.A2(n_1479),
.B1(n_1553),
.B2(n_1594),
.C(n_1617),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1702),
.B(n_1488),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1639),
.B(n_1481),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1639),
.B(n_1481),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1654),
.A2(n_1569),
.B(n_1587),
.C(n_1564),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1633),
.B(n_1601),
.Y(n_1742)
);

BUFx4f_ASAP7_75t_SL g1743 ( 
.A(n_1707),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1631),
.A2(n_1623),
.B(n_1657),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1654),
.A2(n_1577),
.B1(n_1588),
.B2(n_1587),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1722),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1656),
.A2(n_1643),
.B(n_1673),
.C(n_1638),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1646),
.B(n_1469),
.Y(n_1748)
);

AOI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1703),
.A2(n_1588),
.B(n_1569),
.C(n_1483),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1711),
.A2(n_1485),
.B(n_1563),
.C(n_1501),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1722),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1664),
.B(n_1485),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1646),
.B(n_1497),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1635),
.B(n_1574),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1637),
.B(n_1597),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1643),
.A2(n_1551),
.B(n_1568),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1696),
.B(n_1593),
.C(n_1552),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1672),
.B(n_1480),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1664),
.B(n_1582),
.Y(n_1759)
);

AO32x2_ASAP7_75t_L g1760 ( 
.A1(n_1624),
.A2(n_1584),
.A3(n_1632),
.B1(n_1682),
.B2(n_1701),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1637),
.B(n_1647),
.Y(n_1761)
);

BUFx12f_ASAP7_75t_L g1762 ( 
.A(n_1704),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1711),
.A2(n_1684),
.B1(n_1638),
.B2(n_1713),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1703),
.A2(n_1712),
.B(n_1675),
.C(n_1698),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1631),
.A2(n_1641),
.B(n_1657),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1648),
.B(n_1649),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1722),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_L g1768 ( 
.A(n_1722),
.B(n_1671),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_SL g1769 ( 
.A1(n_1732),
.A2(n_1682),
.B(n_1701),
.C(n_1687),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1696),
.A2(n_1698),
.B(n_1685),
.C(n_1687),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1655),
.A2(n_1694),
.B1(n_1693),
.B2(n_1675),
.C(n_1659),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1645),
.B(n_1630),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1712),
.A2(n_1710),
.B1(n_1695),
.B2(n_1705),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1650),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1710),
.A2(n_1705),
.B1(n_1655),
.B2(n_1714),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1713),
.A2(n_1714),
.B(n_1668),
.C(n_1706),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1660),
.B(n_1659),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1685),
.B(n_1627),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1627),
.B(n_1644),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1644),
.B(n_1693),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1658),
.B(n_1726),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1694),
.B(n_1674),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1674),
.B(n_1629),
.Y(n_1783)
);

AOI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1709),
.A2(n_1666),
.B(n_1728),
.Y(n_1784)
);

BUFx2_ASAP7_75t_R g1785 ( 
.A(n_1658),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1700),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1652),
.B(n_1653),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1706),
.A2(n_1699),
.B(n_1671),
.C(n_1680),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1653),
.B(n_1634),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1683),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1699),
.A2(n_1678),
.B(n_1681),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1699),
.A2(n_1697),
.B(n_1671),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1634),
.B(n_1625),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1663),
.B(n_1677),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1678),
.B(n_1681),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1680),
.A2(n_1697),
.B1(n_1724),
.B2(n_1730),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1661),
.B(n_1689),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1708),
.A2(n_1692),
.B(n_1665),
.C(n_1690),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1715),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1717),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1661),
.B(n_1692),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1665),
.B(n_1618),
.Y(n_1803)
);

OA21x2_ASAP7_75t_L g1804 ( 
.A1(n_1628),
.A2(n_1636),
.B(n_1708),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1777),
.B(n_1665),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1787),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1734),
.B(n_1665),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1760),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1783),
.B(n_1665),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1786),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1779),
.B(n_1632),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1783),
.B(n_1642),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1759),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1804),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1782),
.B(n_1642),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1800),
.Y(n_1816)
);

BUFx2_ASAP7_75t_SL g1817 ( 
.A(n_1759),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1779),
.B(n_1768),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1736),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1761),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1743),
.B(n_1704),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1733),
.A2(n_1686),
.B1(n_1688),
.B2(n_1718),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1735),
.B(n_1676),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1804),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1804),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1739),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1798),
.B(n_1802),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1801),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1766),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1802),
.B(n_1716),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1747),
.A2(n_1697),
.B1(n_1680),
.B2(n_1730),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1763),
.A2(n_1686),
.B1(n_1620),
.B2(n_1622),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1795),
.B(n_1679),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1759),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1760),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1764),
.A2(n_1697),
.B1(n_1730),
.B2(n_1719),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1740),
.B(n_1789),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1773),
.A2(n_1725),
.B1(n_1720),
.B2(n_1729),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1790),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1803),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1778),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1746),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1780),
.B(n_1662),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1780),
.B(n_1716),
.Y(n_1845)
);

OAI31xp33_ASAP7_75t_L g1846 ( 
.A1(n_1837),
.A2(n_1750),
.A3(n_1770),
.B(n_1776),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1819),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_SL g1848 ( 
.A(n_1822),
.B(n_1669),
.C(n_1756),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1829),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1809),
.B(n_1751),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1823),
.A2(n_1775),
.B1(n_1791),
.B2(n_1771),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1819),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1818),
.B(n_1811),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1837),
.B(n_1750),
.C(n_1788),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1820),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1814),
.A2(n_1776),
.B(n_1791),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1817),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1809),
.B(n_1767),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1816),
.Y(n_1859)
);

AOI322xp5_ASAP7_75t_L g1860 ( 
.A1(n_1807),
.A2(n_1836),
.A3(n_1808),
.B1(n_1833),
.B2(n_1841),
.C1(n_1781),
.C2(n_1737),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1808),
.B(n_1744),
.C(n_1749),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1810),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1832),
.A2(n_1741),
.B(n_1745),
.C(n_1769),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1814),
.Y(n_1864)
);

NAND4xp25_ASAP7_75t_L g1865 ( 
.A(n_1836),
.B(n_1754),
.C(n_1755),
.D(n_1742),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1818),
.B(n_1767),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_1753),
.Y(n_1867)
);

OAI31xp33_ASAP7_75t_L g1868 ( 
.A1(n_1832),
.A2(n_1799),
.A3(n_1757),
.B(n_1792),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1805),
.B(n_1791),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1814),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1818),
.B(n_1784),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1820),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1829),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1828),
.B(n_1753),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1841),
.B(n_1772),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1825),
.Y(n_1876)
);

INVx4_ASAP7_75t_L g1877 ( 
.A(n_1813),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1843),
.B(n_1744),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1828),
.B(n_1748),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1828),
.B(n_1811),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1840),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1825),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1818),
.B(n_1811),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1845),
.Y(n_1884)
);

BUFx2_ASAP7_75t_L g1885 ( 
.A(n_1811),
.Y(n_1885)
);

AO21x2_ASAP7_75t_L g1886 ( 
.A1(n_1825),
.A2(n_1799),
.B(n_1765),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1840),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1826),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1806),
.Y(n_1889)
);

OAI33xp33_ASAP7_75t_L g1890 ( 
.A1(n_1834),
.A2(n_1796),
.A3(n_1758),
.B1(n_1723),
.B2(n_1721),
.B3(n_1797),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1831),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1839),
.B(n_1744),
.C(n_1754),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1827),
.B(n_1755),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1824),
.B(n_1796),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1838),
.B(n_1794),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1806),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1849),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1847),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1850),
.B(n_1842),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1864),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1846),
.B(n_1835),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1853),
.B(n_1883),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1853),
.B(n_1883),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1861),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1847),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1850),
.B(n_1842),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1849),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1866),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1883),
.B(n_1812),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1883),
.B(n_1844),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1852),
.B(n_1855),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1891),
.B(n_1821),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1873),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1871),
.B(n_1844),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1865),
.B(n_1762),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1872),
.Y(n_1918)
);

AND2x4_ASAP7_75t_SL g1919 ( 
.A(n_1880),
.B(n_1752),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1862),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1881),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1864),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1887),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1884),
.B(n_1830),
.Y(n_1924)
);

INVxp67_ASAP7_75t_SL g1925 ( 
.A(n_1878),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1871),
.B(n_1815),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1887),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1864),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1860),
.B(n_1839),
.C(n_1769),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1896),
.B(n_1830),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1906),
.B(n_1894),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1934)
);

OAI21xp33_ASAP7_75t_L g1935 ( 
.A1(n_1906),
.A2(n_1860),
.B(n_1892),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1900),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1911),
.B(n_1877),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1898),
.B(n_1859),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1900),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1898),
.B(n_1896),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1911),
.B(n_1879),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1917),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1901),
.B(n_1894),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1920),
.B(n_1897),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1907),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1917),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1909),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1909),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1920),
.B(n_1897),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1911),
.B(n_1905),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1905),
.B(n_1879),
.Y(n_1951)
);

INVxp67_ASAP7_75t_L g1952 ( 
.A(n_1915),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1905),
.B(n_1867),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1901),
.B(n_1875),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1907),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1902),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1915),
.B(n_1858),
.Y(n_1957)
);

NOR2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1929),
.B(n_1762),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1925),
.B(n_1918),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1902),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1925),
.B(n_1858),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1903),
.B(n_1893),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1903),
.B(n_1893),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1905),
.B(n_1871),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1913),
.Y(n_1965)
);

INVx2_ASAP7_75t_SL g1966 ( 
.A(n_1919),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1907),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1905),
.B(n_1867),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1919),
.B(n_1874),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1919),
.B(n_1874),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1921),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1918),
.B(n_1889),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1921),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1921),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1923),
.B(n_1889),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1919),
.B(n_1895),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1945),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1952),
.B(n_1930),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1947),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1958),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1944),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1944),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1935),
.A2(n_1929),
.B1(n_1854),
.B2(n_1892),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1945),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1950),
.B(n_1926),
.Y(n_1985)
);

OR2x6_ASAP7_75t_L g1986 ( 
.A(n_1958),
.B(n_1854),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1955),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1948),
.B(n_1930),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1935),
.B(n_1930),
.Y(n_1989)
);

NAND2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1966),
.B(n_1731),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1964),
.B(n_1861),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1938),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1932),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1932),
.B(n_1924),
.Y(n_1994)
);

INVxp67_ASAP7_75t_SL g1995 ( 
.A(n_1942),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1962),
.A2(n_1863),
.B1(n_1851),
.B2(n_1910),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1943),
.B(n_1901),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1950),
.B(n_1926),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1943),
.B(n_1908),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1955),
.Y(n_2000)
);

AND3x2_ASAP7_75t_L g2001 ( 
.A(n_1946),
.B(n_1846),
.C(n_1863),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1963),
.B(n_1865),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1969),
.B(n_1926),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1967),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1966),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1969),
.B(n_1926),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1949),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1949),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1965),
.B(n_1924),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1956),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1940),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1965),
.B(n_1924),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1957),
.B(n_1914),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1983),
.B(n_1954),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_2001),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1995),
.B(n_1954),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1989),
.B(n_1848),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1993),
.B(n_1959),
.Y(n_2018)
);

AOI32xp33_ASAP7_75t_SL g2019 ( 
.A1(n_1980),
.A2(n_1939),
.A3(n_1936),
.B1(n_1959),
.B2(n_1973),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1977),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1979),
.B(n_1964),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_2005),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1977),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1986),
.B(n_1939),
.C(n_1936),
.Y(n_2024)
);

NOR3xp33_ASAP7_75t_L g2025 ( 
.A(n_1991),
.B(n_1961),
.C(n_1890),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1986),
.A2(n_1868),
.B(n_1890),
.Y(n_2026)
);

AOI21xp33_ASAP7_75t_SL g2027 ( 
.A1(n_1986),
.A2(n_1910),
.B(n_1964),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1992),
.B(n_1941),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1984),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_2005),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1984),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1986),
.B(n_1953),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_2008),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_2010),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1985),
.B(n_1953),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1996),
.A2(n_1878),
.B1(n_1869),
.B2(n_1956),
.C(n_1960),
.Y(n_2036)
);

OAI32xp33_ASAP7_75t_L g2037 ( 
.A1(n_2002),
.A2(n_1971),
.A3(n_1967),
.B1(n_1974),
.B2(n_1973),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1978),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1987),
.Y(n_2039)
);

INVxp33_ASAP7_75t_L g2040 ( 
.A(n_1988),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2011),
.B(n_1941),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1997),
.B(n_1972),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2026),
.A2(n_2014),
.B1(n_2025),
.B2(n_2024),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2020),
.Y(n_2044)
);

O2A1O1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_2037),
.A2(n_1981),
.B(n_2007),
.C(n_1982),
.Y(n_2045)
);

NAND2x1_ASAP7_75t_L g2046 ( 
.A(n_2035),
.B(n_1985),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2020),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2031),
.Y(n_2048)
);

OAI21xp33_ASAP7_75t_L g2049 ( 
.A1(n_2032),
.A2(n_1994),
.B(n_2009),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2030),
.B(n_1997),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2035),
.B(n_1998),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_2040),
.A2(n_1999),
.B1(n_1998),
.B2(n_1910),
.Y(n_2052)
);

OAI22xp33_ASAP7_75t_SL g2053 ( 
.A1(n_2015),
.A2(n_2018),
.B1(n_2016),
.B2(n_2021),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_SL g2054 ( 
.A(n_2036),
.B(n_2015),
.C(n_2027),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2022),
.B(n_1999),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2017),
.A2(n_2034),
.B1(n_2028),
.B2(n_2041),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2031),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2039),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2039),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2037),
.A2(n_2012),
.B(n_1868),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_2018),
.B(n_2013),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2033),
.A2(n_2006),
.B1(n_2003),
.B2(n_1970),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2023),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2017),
.B(n_2004),
.C(n_2000),
.D(n_1987),
.Y(n_2064)
);

XNOR2xp5_ASAP7_75t_L g2065 ( 
.A(n_2043),
.B(n_2038),
.Y(n_2065)
);

OAI21xp33_ASAP7_75t_L g2066 ( 
.A1(n_2060),
.A2(n_2042),
.B(n_2006),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2046),
.Y(n_2067)
);

AOI322xp5_ASAP7_75t_L g2068 ( 
.A1(n_2054),
.A2(n_2019),
.A3(n_2034),
.B1(n_2010),
.B2(n_2029),
.C1(n_1960),
.C2(n_1956),
.Y(n_2068)
);

AOI322xp5_ASAP7_75t_L g2069 ( 
.A1(n_2061),
.A2(n_2019),
.A3(n_1960),
.B1(n_1869),
.B2(n_2000),
.C1(n_2004),
.C2(n_1870),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2055),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2050),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2044),
.Y(n_2072)
);

NAND2x1_ASAP7_75t_L g2073 ( 
.A(n_2051),
.B(n_2003),
.Y(n_2073)
);

OAI21xp33_ASAP7_75t_L g2074 ( 
.A1(n_2053),
.A2(n_2042),
.B(n_1964),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2047),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2048),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2057),
.Y(n_2077)
);

OAI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2064),
.A2(n_1990),
.B(n_1974),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2074),
.A2(n_2045),
.B1(n_2064),
.B2(n_2049),
.C(n_2056),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_2071),
.A2(n_2059),
.B(n_2058),
.C(n_2063),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2077),
.Y(n_2081)
);

AOI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2066),
.A2(n_2052),
.B1(n_2062),
.B2(n_1971),
.C(n_1871),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2073),
.B(n_1968),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_2067),
.Y(n_2084)
);

AOI211xp5_ASAP7_75t_L g2085 ( 
.A1(n_2065),
.A2(n_1738),
.B(n_1916),
.C(n_1970),
.Y(n_2085)
);

NAND3xp33_ASAP7_75t_L g2086 ( 
.A(n_2068),
.B(n_1933),
.C(n_1931),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2077),
.A2(n_1856),
.B1(n_1886),
.B2(n_1902),
.Y(n_2087)
);

NOR2xp67_ASAP7_75t_L g2088 ( 
.A(n_2070),
.B(n_1968),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_2069),
.B(n_1990),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_2081),
.B(n_2072),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2079),
.A2(n_2078),
.B(n_2076),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2089),
.A2(n_2078),
.B(n_2075),
.Y(n_2092)
);

AOI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_2080),
.A2(n_1870),
.B1(n_1928),
.B2(n_1902),
.C(n_1922),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2083),
.Y(n_2094)
);

A2O1A1Ixp33_ASAP7_75t_L g2095 ( 
.A1(n_2088),
.A2(n_1928),
.B(n_1922),
.C(n_1785),
.Y(n_2095)
);

AOI221xp5_ASAP7_75t_L g2096 ( 
.A1(n_2086),
.A2(n_1922),
.B1(n_1928),
.B2(n_1990),
.C(n_1856),
.Y(n_2096)
);

AOI211xp5_ASAP7_75t_L g2097 ( 
.A1(n_2091),
.A2(n_2092),
.B(n_2084),
.C(n_2095),
.Y(n_2097)
);

AOI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2094),
.A2(n_2082),
.B(n_2085),
.C(n_1916),
.Y(n_2098)
);

AOI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_2096),
.A2(n_2087),
.B1(n_1928),
.B2(n_1922),
.C(n_1856),
.Y(n_2099)
);

AOI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2093),
.A2(n_1856),
.B1(n_1975),
.B2(n_1972),
.C(n_1882),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2090),
.A2(n_1975),
.B(n_1933),
.Y(n_2101)
);

AOI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2092),
.A2(n_1876),
.B1(n_1882),
.B2(n_1888),
.C(n_1886),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2090),
.Y(n_2103)
);

AOI221xp5_ASAP7_75t_L g2104 ( 
.A1(n_2092),
.A2(n_1876),
.B1(n_1882),
.B2(n_1888),
.C(n_1886),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2103),
.B(n_1951),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2101),
.B(n_1951),
.Y(n_2106)
);

AND2x2_ASAP7_75t_SL g2107 ( 
.A(n_2097),
.B(n_1731),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2098),
.Y(n_2108)
);

AO22x1_ASAP7_75t_L g2109 ( 
.A1(n_2102),
.A2(n_1934),
.B1(n_1931),
.B2(n_1937),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2104),
.A2(n_1916),
.B1(n_1857),
.B2(n_1926),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_2107),
.B(n_2099),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_L g2112 ( 
.A(n_2108),
.B(n_2100),
.C(n_1934),
.Y(n_2112)
);

OR4x1_ASAP7_75t_L g2113 ( 
.A(n_2105),
.B(n_1923),
.C(n_1927),
.D(n_1937),
.Y(n_2113)
);

CKINVDCx16_ASAP7_75t_R g2114 ( 
.A(n_2113),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_2114),
.Y(n_2115)
);

OAI22x1_ASAP7_75t_L g2116 ( 
.A1(n_2115),
.A2(n_2112),
.B1(n_2111),
.B2(n_2106),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2115),
.A2(n_2110),
.B1(n_2109),
.B2(n_1908),
.Y(n_2117)
);

OAI22x1_ASAP7_75t_L g2118 ( 
.A1(n_2116),
.A2(n_1916),
.B1(n_1976),
.B2(n_1724),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2117),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2118),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2119),
.B(n_1899),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2121),
.B(n_1916),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2122),
.B(n_2120),
.Y(n_2123)
);

NAND3x2_ASAP7_75t_L g2124 ( 
.A(n_2123),
.B(n_1899),
.C(n_1976),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_R g2125 ( 
.A1(n_2124),
.A2(n_1899),
.B1(n_1817),
.B2(n_1908),
.C(n_1912),
.Y(n_2125)
);

AOI211xp5_ASAP7_75t_L g2126 ( 
.A1(n_2125),
.A2(n_1730),
.B(n_1729),
.C(n_1727),
.Y(n_2126)
);


endmodule