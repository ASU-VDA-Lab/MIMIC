module fake_aes_7697_n_1436 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1436);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1436;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1130;
wire n_584;
wire n_1042;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVxp67_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_116), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_37), .Y(n_306) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_242), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_213), .B(n_232), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_191), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_170), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_167), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_109), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_78), .Y(n_314) );
CKINVDCx14_ASAP7_75t_R g315 ( .A(n_252), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_214), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_276), .Y(n_317) );
INVxp33_ASAP7_75t_L g318 ( .A(n_152), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_96), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_38), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_212), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_196), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_187), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_74), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_39), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_221), .B(n_96), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_80), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_203), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_302), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_95), .Y(n_330) );
INVxp33_ASAP7_75t_L g331 ( .A(n_193), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_231), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_35), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_88), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_6), .Y(n_335) );
INVxp33_ASAP7_75t_SL g336 ( .A(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_148), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_178), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_299), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_63), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_48), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_223), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_154), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_184), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_274), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_26), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_62), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_37), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_124), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_150), .B(n_257), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_160), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_281), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_43), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_50), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_45), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_22), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_180), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_79), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_198), .Y(n_359) );
INVxp33_ASAP7_75t_SL g360 ( .A(n_296), .Y(n_360) );
INVxp33_ASAP7_75t_L g361 ( .A(n_179), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_279), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_175), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_205), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_77), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_92), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_95), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_18), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_88), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_247), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_108), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_173), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_256), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_201), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_56), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_3), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_225), .Y(n_377) );
INVxp33_ASAP7_75t_L g378 ( .A(n_216), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_28), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_9), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_27), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_8), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_113), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_222), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_66), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_6), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_137), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_224), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_65), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_215), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_123), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_103), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_46), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_55), .Y(n_394) );
CKINVDCx14_ASAP7_75t_R g395 ( .A(n_7), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_192), .B(n_99), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_42), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_163), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_112), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_71), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_10), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_235), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_22), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_8), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_86), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_33), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_49), .Y(n_407) );
INVxp33_ASAP7_75t_L g408 ( .A(n_195), .Y(n_408) );
INVxp33_ASAP7_75t_SL g409 ( .A(n_141), .Y(n_409) );
INVxp33_ASAP7_75t_L g410 ( .A(n_86), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_136), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_82), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_135), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_0), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_258), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_93), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_42), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_140), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_261), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_5), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_298), .Y(n_421) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_61), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_66), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_219), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_218), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_107), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_69), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_146), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_145), .Y(n_429) );
INVxp33_ASAP7_75t_L g430 ( .A(n_44), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_204), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_185), .B(n_275), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_144), .Y(n_433) );
INVxp33_ASAP7_75t_SL g434 ( .A(n_85), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_84), .Y(n_435) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_206), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_67), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_271), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_149), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_228), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_100), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_110), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_292), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_7), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_283), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_220), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_5), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_106), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_19), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_71), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_139), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_169), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_419), .Y(n_454) );
NAND2xp33_ASAP7_75t_R g455 ( .A(n_336), .B(n_0), .Y(n_455) );
NOR2xp33_ASAP7_75t_R g456 ( .A(n_315), .B(n_97), .Y(n_456) );
AND2x6_ASAP7_75t_L g457 ( .A(n_313), .B(n_98), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_395), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_334), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_334), .B(n_1), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_407), .B(n_1), .Y(n_462) );
NOR2xp67_ASAP7_75t_L g463 ( .A(n_363), .B(n_2), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_373), .B(n_2), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_411), .B(n_3), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_349), .Y(n_466) );
NOR2xp33_ASAP7_75t_SL g467 ( .A(n_445), .B(n_316), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_309), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_309), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_410), .B(n_4), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_314), .B(n_4), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_311), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_326), .B(n_101), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_311), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_369), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_9), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_374), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_433), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_419), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_314), .B(n_10), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_312), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_316), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_312), .Y(n_484) );
NOR2xp33_ASAP7_75t_SL g485 ( .A(n_321), .B(n_301), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_436), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_419), .Y(n_487) );
INVx4_ASAP7_75t_SL g488 ( .A(n_457), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_458), .B(n_330), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_457), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_460), .B(n_330), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_480), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_486), .B(n_321), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_458), .B(n_304), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_453), .B(n_461), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_483), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
INVx4_ASAP7_75t_SL g501 ( .A(n_457), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_486), .B(n_332), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_480), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_476), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_460), .B(n_318), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_461), .B(n_319), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_476), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_476), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_470), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_467), .B(n_332), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_461), .B(n_447), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_480), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_468), .B(n_319), .Y(n_514) );
BUFx3_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_480), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_468), .B(n_304), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_476), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
AO22x2_ASAP7_75t_L g522 ( .A1(n_469), .A2(n_322), .B1(n_323), .B2(n_317), .Y(n_522) );
AO22x2_ASAP7_75t_L g523 ( .A1(n_469), .A2(n_322), .B1(n_323), .B2(n_317), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g525 ( .A1(n_466), .A2(n_397), .B1(n_434), .B2(n_325), .Y(n_525) );
AND2x6_ASAP7_75t_L g526 ( .A(n_470), .B(n_326), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_487), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_470), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_477), .B(n_331), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_472), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_487), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_477), .B(n_361), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_490), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_499), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_512), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_488), .B(n_474), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_488), .B(n_474), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g541 ( .A(n_525), .B(n_479), .C(n_478), .Y(n_541) );
INVx8_ASAP7_75t_L g542 ( .A(n_526), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_490), .Y(n_543) );
AND3x1_ASAP7_75t_SL g544 ( .A(n_525), .B(n_367), .C(n_365), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_526), .Y(n_545) );
OR2x2_ASAP7_75t_SL g546 ( .A(n_509), .B(n_354), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_526), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_489), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_488), .B(n_474), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_498), .B(n_477), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_526), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_526), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_498), .B(n_463), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_526), .A2(n_455), .B1(n_459), .B2(n_464), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_490), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_499), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_522), .A2(n_482), .B1(n_484), .B2(n_475), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_509), .A2(n_465), .B(n_464), .C(n_471), .Y(n_561) );
NOR3xp33_ASAP7_75t_SL g562 ( .A(n_495), .B(n_455), .C(n_450), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_491), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_498), .B(n_475), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_526), .Y(n_565) );
INVx4_ASAP7_75t_L g566 ( .A(n_526), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_494), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_498), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
NOR2xp33_ASAP7_75t_R g570 ( .A(n_526), .B(n_459), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_498), .B(n_482), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_500), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_497), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_512), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_505), .B(n_484), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_505), .B(n_534), .Y(n_579) );
INVxp33_ASAP7_75t_L g580 ( .A(n_512), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_491), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_506), .B(n_463), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_531), .B(n_465), .Y(n_583) );
BUFx10_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_506), .B(n_471), .Y(n_586) );
INVx6_ASAP7_75t_L g587 ( .A(n_514), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_534), .B(n_462), .Y(n_588) );
AND3x1_ASAP7_75t_SL g589 ( .A(n_492), .B(n_379), .C(n_375), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_529), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_514), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_514), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_514), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_522), .Y(n_595) );
NOR3xp33_ASAP7_75t_SL g596 ( .A(n_502), .B(n_355), .C(n_348), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_506), .B(n_481), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_522), .Y(n_599) );
AND3x1_ASAP7_75t_SL g600 ( .A(n_492), .B(n_381), .C(n_380), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_515), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_531), .B(n_348), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_531), .B(n_462), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_515), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_530), .A2(n_474), .B(n_432), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_534), .B(n_481), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_521), .Y(n_607) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_532), .Y(n_608) );
NAND2xp33_ASAP7_75t_SL g609 ( .A(n_532), .B(n_456), .Y(n_609) );
BUFx8_ASAP7_75t_L g610 ( .A(n_492), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_506), .B(n_344), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_522), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_521), .A2(n_434), .B1(n_355), .B2(n_485), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_510), .B(n_378), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_496), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_518), .B(n_366), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_518), .B(n_408), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_496), .B(n_344), .Y(n_619) );
OR2x6_ASAP7_75t_L g620 ( .A(n_523), .B(n_335), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_523), .B(n_371), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_523), .B(n_371), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_523), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_507), .B(n_306), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_507), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_605), .A2(n_515), .B(n_523), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_537), .B(n_590), .Y(n_628) );
INVx3_ASAP7_75t_SL g629 ( .A(n_559), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_542), .Y(n_630) );
BUFx10_ASAP7_75t_L g631 ( .A(n_559), .Y(n_631) );
BUFx8_ASAP7_75t_L g632 ( .A(n_556), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_543), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_566), .B(n_488), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_591), .A2(n_485), .B1(n_336), .B2(n_409), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_610), .Y(n_637) );
BUFx3_ASAP7_75t_L g638 ( .A(n_610), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_539), .A2(n_508), .B(n_504), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_612), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_566), .Y(n_641) );
INVx4_ASAP7_75t_L g642 ( .A(n_542), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_616), .B(n_360), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_591), .Y(n_644) );
BUFx12f_ASAP7_75t_L g645 ( .A(n_610), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_566), .B(n_396), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx5_ASAP7_75t_L g648 ( .A(n_542), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_543), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_570), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_620), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_583), .B(n_333), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_542), .Y(n_653) );
OR2x6_ASAP7_75t_L g654 ( .A(n_545), .B(n_320), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_617), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_543), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_541), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_579), .B(n_360), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_539), .A2(n_508), .B(n_504), .Y(n_659) );
BUFx12f_ASAP7_75t_L g660 ( .A(n_546), .Y(n_660) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_601), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_586), .B(n_409), .Y(n_662) );
BUFx12f_ASAP7_75t_L g663 ( .A(n_582), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_584), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_585), .A2(n_528), .B(n_519), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_587), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_562), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_584), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_585), .A2(n_528), .B(n_519), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_549), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_570), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_576), .B(n_403), .Y(n_672) );
BUFx4f_ASAP7_75t_L g673 ( .A(n_620), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_540), .A2(n_308), .B(n_328), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_620), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_545), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_538), .A2(n_420), .B1(n_422), .B2(n_376), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_555), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_602), .B(n_320), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_586), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_587), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_580), .B(n_324), .Y(n_684) );
INVx4_ASAP7_75t_L g685 ( .A(n_555), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_565), .Y(n_686) );
INVxp67_ASAP7_75t_L g687 ( .A(n_586), .Y(n_687) );
INVx4_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_598), .B(n_456), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_598), .B(n_425), .Y(n_690) );
INVx8_ASAP7_75t_L g691 ( .A(n_598), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_560), .B(n_488), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_548), .B(n_396), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_596), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_588), .B(n_425), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_606), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_603), .B(n_385), .Y(n_697) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_563), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_563), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_549), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_550), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_535), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_607), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_618), .B(n_389), .Y(n_704) );
OR2x6_ASAP7_75t_L g705 ( .A(n_554), .B(n_324), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_560), .B(n_488), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_580), .B(n_340), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_624), .Y(n_708) );
INVx5_ASAP7_75t_L g709 ( .A(n_568), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_582), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g711 ( .A1(n_553), .A2(n_406), .B1(n_449), .B2(n_444), .C1(n_437), .C2(n_358), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_536), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_595), .A2(n_457), .B1(n_341), .B2(n_346), .Y(n_713) );
BUFx2_ASAP7_75t_R g714 ( .A(n_607), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_556), .B(n_501), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_547), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_563), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_582), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_609), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_557), .A2(n_394), .B1(n_400), .B2(n_393), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_558), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_611), .B(n_340), .Y(n_722) );
BUFx4f_ASAP7_75t_L g723 ( .A(n_556), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_568), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_614), .Y(n_725) );
INVx4_ASAP7_75t_L g726 ( .A(n_569), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_618), .A2(n_412), .B1(n_414), .B2(n_401), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_578), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_615), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_592), .Y(n_730) );
INVx1_ASAP7_75t_SL g731 ( .A(n_625), .Y(n_731) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_597), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_577), .B(n_341), .Y(n_733) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_569), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_599), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_561), .B(n_435), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_613), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_622), .A2(n_594), .B1(n_593), .B2(n_572), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_540), .A2(n_329), .B(n_328), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_564), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_551), .A2(n_337), .B(n_329), .Y(n_741) );
AOI21x1_ASAP7_75t_L g742 ( .A1(n_551), .A2(n_511), .B(n_503), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_619), .B(n_346), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_608), .B(n_347), .Y(n_744) );
AO21x1_ASAP7_75t_L g745 ( .A1(n_621), .A2(n_338), .B(n_337), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_609), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_623), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_550), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_615), .B(n_347), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_552), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_569), .Y(n_751) );
BUFx8_ASAP7_75t_L g752 ( .A(n_544), .Y(n_752) );
AO22x2_ASAP7_75t_L g753 ( .A1(n_589), .A2(n_356), .B1(n_358), .B2(n_353), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_573), .A2(n_457), .B1(n_356), .B2(n_368), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_574), .A2(n_339), .B(n_338), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_552), .B(n_501), .Y(n_756) );
CKINVDCx12_ASAP7_75t_R g757 ( .A(n_600), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_567), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_567), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_569), .Y(n_760) );
AO21x1_ASAP7_75t_L g761 ( .A1(n_571), .A2(n_343), .B(n_339), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g762 ( .A1(n_711), .A2(n_353), .B(n_404), .C(n_368), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_696), .B(n_571), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_648), .B(n_575), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_670), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_700), .Y(n_766) );
CKINVDCx11_ASAP7_75t_R g767 ( .A(n_629), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_SL g768 ( .A1(n_658), .A2(n_350), .B(n_575), .C(n_507), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_645), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_753), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_673), .A2(n_404), .B1(n_416), .B2(n_406), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_753), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_655), .A2(n_437), .B1(n_444), .B2(n_423), .C(n_416), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_673), .A2(n_369), .B1(n_449), .B2(n_423), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_740), .A2(n_369), .B1(n_382), .B2(n_327), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_SL g776 ( .A1(n_750), .A2(n_305), .B(n_372), .C(n_364), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_627), .A2(n_626), .B(n_457), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_740), .B(n_626), .Y(n_778) );
INVx6_ASAP7_75t_L g779 ( .A(n_632), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_628), .B(n_327), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_644), .B(n_382), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_629), .B(n_386), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_753), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_744), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_637), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_703), .A2(n_369), .B1(n_405), .B2(n_386), .Y(n_786) );
BUFx12f_ASAP7_75t_L g787 ( .A(n_631), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_658), .A2(n_369), .B1(n_417), .B2(n_405), .Y(n_788) );
O2A1O1Ixp5_ASAP7_75t_L g789 ( .A1(n_745), .A2(n_359), .B(n_473), .C(n_454), .Y(n_789) );
INVx4_ASAP7_75t_L g790 ( .A(n_691), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_701), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_748), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_758), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_747), .A2(n_427), .B1(n_417), .B2(n_457), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_684), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_731), .B(n_427), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_649), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_691), .B(n_581), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_691), .B(n_581), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_680), .A2(n_457), .B1(n_343), .B2(n_352), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_652), .A2(n_303), .B1(n_415), .B2(n_421), .C(n_443), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_680), .A2(n_604), .B1(n_581), .B2(n_310), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_631), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_637), .Y(n_804) );
INVxp33_ASAP7_75t_L g805 ( .A(n_672), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_707), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g807 ( .A1(n_679), .A2(n_421), .B1(n_448), .B2(n_345), .C(n_443), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_687), .A2(n_457), .B1(n_352), .B2(n_357), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_703), .A2(n_313), .B1(n_398), .B2(n_383), .Y(n_809) );
CKINVDCx6p67_ASAP7_75t_R g810 ( .A(n_638), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_643), .B(n_11), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_729), .B(n_581), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_702), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_687), .B(n_604), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_657), .Y(n_815) );
NAND2xp33_ASAP7_75t_R g816 ( .A(n_651), .B(n_11), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_712), .Y(n_817) );
INVx2_ASAP7_75t_SL g818 ( .A(n_632), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_675), .A2(n_398), .B1(n_442), .B2(n_383), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_704), .A2(n_415), .B1(n_452), .B2(n_345), .C(n_446), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g821 ( .A1(n_705), .A2(n_362), .B1(n_402), .B2(n_357), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_716), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_649), .Y(n_823) );
INVx2_ASAP7_75t_SL g824 ( .A(n_663), .Y(n_824) );
NAND2x1p5_ASAP7_75t_L g825 ( .A(n_648), .B(n_604), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_695), .B(n_12), .Y(n_826) );
INVx2_ASAP7_75t_SL g827 ( .A(n_723), .Y(n_827) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_750), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_733), .B(n_12), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_759), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_727), .A2(n_307), .B1(n_342), .B2(n_351), .C(n_438), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_705), .B(n_13), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_738), .A2(n_362), .B1(n_424), .B2(n_402), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_721), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_705), .A2(n_439), .B1(n_440), .B2(n_424), .Y(n_835) );
INVx4_ASAP7_75t_L g836 ( .A(n_648), .Y(n_836) );
A2O1A1Ixp33_ASAP7_75t_L g837 ( .A1(n_739), .A2(n_440), .B(n_441), .C(n_439), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_648), .B(n_501), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_738), .A2(n_446), .B1(n_448), .B2(n_441), .Y(n_839) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_654), .B(n_452), .Y(n_840) );
BUFx3_ASAP7_75t_L g841 ( .A(n_660), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_752), .A2(n_442), .B1(n_370), .B2(n_384), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_735), .A2(n_377), .B1(n_388), .B2(n_387), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_714), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_654), .A2(n_390), .B1(n_392), .B2(n_391), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_728), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_662), .B(n_604), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_720), .B(n_399), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_752), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_634), .Y(n_850) );
INVxp67_ASAP7_75t_L g851 ( .A(n_708), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g852 ( .A(n_709), .B(n_501), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_627), .A2(n_501), .B(n_503), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_646), .A2(n_413), .B1(n_426), .B2(n_418), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_730), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_749), .B(n_428), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_654), .Y(n_857) );
OAI21x1_ASAP7_75t_L g858 ( .A1(n_742), .A2(n_359), .B(n_429), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_642), .B(n_501), .Y(n_859) );
CKINVDCx16_ASAP7_75t_R g860 ( .A(n_650), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_640), .A2(n_431), .B1(n_451), .B2(n_419), .Y(n_861) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_739), .A2(n_507), .B(n_473), .C(n_454), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_722), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_761), .A2(n_473), .A3(n_454), .B(n_503), .Y(n_864) );
AO31x2_ASAP7_75t_L g865 ( .A1(n_741), .A2(n_511), .A3(n_517), .B(n_516), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_725), .B(n_13), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_757), .A2(n_507), .B1(n_487), .B2(n_511), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_708), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_736), .Y(n_869) );
CKINVDCx6p67_ASAP7_75t_R g870 ( .A(n_650), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_640), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_681), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_642), .B(n_14), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_656), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_697), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_743), .Y(n_876) );
AOI221xp5_ASAP7_75t_SL g877 ( .A1(n_755), .A2(n_487), .B1(n_527), .B2(n_524), .C(n_517), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_710), .Y(n_878) );
BUFx3_ASAP7_75t_L g879 ( .A(n_647), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_671), .A2(n_487), .B1(n_517), .B2(n_516), .Y(n_880) );
CKINVDCx6p67_ASAP7_75t_R g881 ( .A(n_671), .Y(n_881) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_646), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_667), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_735), .A2(n_737), .B1(n_718), .B2(n_732), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_737), .A2(n_487), .B1(n_524), .B2(n_516), .Y(n_885) );
CKINVDCx11_ASAP7_75t_R g886 ( .A(n_630), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_694), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_724), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_732), .A2(n_487), .B1(n_527), .B2(n_524), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_674), .A2(n_527), .B(n_513), .Y(n_890) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_683), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_690), .B(n_14), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_709), .Y(n_893) );
OAI211xp5_ASAP7_75t_SL g894 ( .A1(n_677), .A2(n_15), .B(n_16), .C(n_17), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_755), .A2(n_487), .B1(n_520), .B2(n_513), .C(n_493), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_723), .B(n_15), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_666), .Y(n_897) );
AND2x6_ASAP7_75t_L g898 ( .A(n_630), .B(n_493), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_751), .Y(n_899) );
OAI22xp33_ASAP7_75t_L g900 ( .A1(n_693), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_693), .B(n_19), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_636), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_639), .A2(n_513), .B(n_493), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_633), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_689), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_751), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_719), .A2(n_533), .B1(n_520), .B2(n_513), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_674), .A2(n_513), .B(n_493), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_770), .A2(n_772), .B1(n_783), .B2(n_894), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_863), .B(n_664), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_813), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_763), .B(n_668), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_830), .Y(n_913) );
INVx3_ASAP7_75t_L g914 ( .A(n_836), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_875), .B(n_746), .Y(n_915) );
BUFx12f_ASAP7_75t_L g916 ( .A(n_767), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_876), .B(n_668), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g918 ( .A1(n_821), .A2(n_653), .B1(n_709), .B2(n_741), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_882), .A2(n_709), .B1(n_692), .B2(n_706), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_882), .A2(n_692), .B1(n_706), .B2(n_653), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_821), .A2(n_713), .B1(n_754), .B2(n_686), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_786), .A2(n_686), .B1(n_676), .B2(n_685), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_786), .A2(n_676), .B1(n_688), .B2(n_685), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_869), .A2(n_902), .B1(n_829), .B2(n_795), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_817), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_790), .B(n_630), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_902), .A2(n_806), .B1(n_784), .B2(n_773), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_805), .B(n_688), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_779), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_866), .B(n_24), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_835), .A2(n_713), .B1(n_754), .B2(n_661), .Y(n_931) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_771), .A2(n_641), .B1(n_669), .B2(n_665), .C(n_678), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_788), .A2(n_678), .B1(n_641), .B2(n_661), .Y(n_933) );
AOI221xp5_ASAP7_75t_SL g934 ( .A1(n_845), .A2(n_639), .B1(n_659), .B2(n_661), .C(n_682), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_789), .A2(n_659), .B(n_756), .Y(n_935) );
INVx4_ASAP7_75t_L g936 ( .A(n_886), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_765), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_828), .B(n_780), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_835), .A2(n_661), .B1(n_682), .B2(n_630), .Y(n_939) );
OAI21xp33_ASAP7_75t_SL g940 ( .A1(n_840), .A2(n_726), .B(n_698), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_790), .B(n_715), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_831), .A2(n_682), .B1(n_715), .B2(n_726), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_828), .A2(n_682), .B1(n_760), .B2(n_734), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_845), .A2(n_635), .B1(n_756), .B2(n_734), .Y(n_944) );
OA21x2_ASAP7_75t_L g945 ( .A1(n_877), .A2(n_635), .B(n_683), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_832), .A2(n_760), .B1(n_734), .B2(n_717), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_873), .A2(n_760), .B1(n_734), .B2(n_717), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_822), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_834), .B(n_760), .Y(n_949) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_900), .A2(n_24), .A3(n_25), .B1(n_26), .B2(n_27), .B3(n_28), .Y(n_950) );
OR2x6_ASAP7_75t_L g951 ( .A(n_779), .B(n_683), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_771), .A2(n_717), .B1(n_699), .B2(n_698), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_873), .A2(n_717), .B1(n_699), .B2(n_698), .Y(n_953) );
BUFx2_ASAP7_75t_L g954 ( .A(n_785), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g955 ( .A1(n_857), .A2(n_699), .B1(n_698), .B2(n_683), .Y(n_955) );
OAI221xp5_ASAP7_75t_SL g956 ( .A1(n_900), .A2(n_25), .B1(n_29), .B2(n_30), .C(n_31), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_766), .Y(n_957) );
OA21x2_ASAP7_75t_L g958 ( .A1(n_903), .A2(n_699), .B(n_513), .Y(n_958) );
INVx4_ASAP7_75t_L g959 ( .A(n_779), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_782), .B(n_29), .Y(n_960) );
OAI21xp33_ASAP7_75t_L g961 ( .A1(n_809), .A2(n_513), .B(n_493), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_791), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_801), .A2(n_533), .B1(n_520), .B2(n_493), .C(n_33), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_871), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_781), .B(n_32), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_836), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_788), .A2(n_533), .B1(n_520), .B2(n_493), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_871), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_816), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_969) );
INVx4_ASAP7_75t_L g970 ( .A(n_769), .Y(n_970) );
NAND3xp33_ASAP7_75t_L g971 ( .A(n_809), .B(n_533), .C(n_520), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_826), .A2(n_533), .B1(n_520), .B2(n_38), .Y(n_972) );
AO31x2_ASAP7_75t_L g973 ( .A1(n_853), .A2(n_34), .A3(n_36), .B(n_39), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_846), .B(n_40), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_842), .A2(n_533), .B1(n_520), .B2(n_43), .C(n_44), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_868), .B(n_40), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_901), .A2(n_533), .B1(n_45), .B2(n_46), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_855), .Y(n_978) );
AOI21xp33_ASAP7_75t_SL g979 ( .A1(n_844), .A2(n_41), .B(n_47), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_854), .A2(n_41), .B1(n_47), .B2(n_48), .Y(n_980) );
AOI222xp33_ASAP7_75t_L g981 ( .A1(n_762), .A2(n_49), .B1(n_50), .B2(n_51), .C1(n_52), .C2(n_53), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_804), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_807), .A2(n_51), .B1(n_52), .B2(n_53), .C(n_54), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_868), .A2(n_811), .B1(n_896), .B2(n_818), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_904), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g986 ( .A1(n_908), .A2(n_104), .B(n_102), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_796), .B(n_54), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_905), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_884), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_989) );
INVx2_ASAP7_75t_SL g990 ( .A(n_787), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_820), .A2(n_892), .B1(n_833), .B2(n_839), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_792), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_851), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_993) );
OAI22xp5_ASAP7_75t_SL g994 ( .A1(n_842), .A2(n_860), .B1(n_849), .B2(n_887), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_872), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_851), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_996) );
AOI222xp33_ASAP7_75t_L g997 ( .A1(n_848), .A2(n_63), .B1(n_64), .B2(n_65), .C1(n_67), .C2(n_68), .Y(n_997) );
OAI21x1_ASAP7_75t_L g998 ( .A1(n_858), .A2(n_111), .B(n_105), .Y(n_998) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_778), .A2(n_64), .B1(n_68), .B2(n_69), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_824), .B(n_70), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_768), .B(n_70), .C(n_72), .Y(n_1001) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_841), .A2(n_72), .B1(n_73), .B2(n_74), .C1(n_75), .C2(n_76), .Y(n_1002) );
INVx3_ASAP7_75t_L g1003 ( .A(n_764), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_893), .A2(n_73), .B1(n_75), .B2(n_76), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_793), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_888), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_803), .B(n_77), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_789), .A2(n_78), .B(n_79), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_833), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_1009) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_856), .A2(n_839), .B1(n_878), .B2(n_883), .C1(n_774), .C2(n_897), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_870), .B(n_81), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_850), .Y(n_1012) );
OAI211xp5_ASAP7_75t_L g1013 ( .A1(n_819), .A2(n_774), .B(n_861), .C(n_775), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_893), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1015 ( .A1(n_867), .A2(n_83), .B1(n_87), .B2(n_89), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_879), .B(n_87), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_812), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_827), .B(n_90), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_874), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_775), .Y(n_1020) );
INVx5_ASAP7_75t_SL g1021 ( .A(n_810), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_884), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_1022) );
INVx3_ASAP7_75t_L g1023 ( .A(n_764), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_881), .B(n_94), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1025 ( .A1(n_837), .A2(n_94), .B(n_114), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_843), .A2(n_115), .B1(n_117), .B2(n_118), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_865), .Y(n_1027) );
OAI22xp33_ASAP7_75t_L g1028 ( .A1(n_777), .A2(n_119), .B1(n_120), .B2(n_121), .Y(n_1028) );
BUFx4f_ASAP7_75t_SL g1029 ( .A(n_898), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_865), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_843), .A2(n_122), .B1(n_125), .B2(n_126), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_815), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_859), .B(n_127), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_819), .B(n_128), .Y(n_1034) );
INVx3_ASAP7_75t_L g1035 ( .A(n_898), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g1036 ( .A1(n_890), .A2(n_776), .B(n_862), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_797), .B(n_129), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_861), .A2(n_130), .B1(n_131), .B2(n_132), .C(n_133), .Y(n_1038) );
AOI221x1_ASAP7_75t_SL g1039 ( .A1(n_847), .A2(n_134), .B1(n_138), .B2(n_142), .C(n_143), .Y(n_1039) );
NAND2xp33_ASAP7_75t_L g1040 ( .A(n_898), .B(n_147), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_823), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_968), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1043 ( .A1(n_927), .A2(n_794), .B(n_800), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_1010), .A2(n_794), .B1(n_802), .B2(n_808), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_968), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_1029), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1027), .Y(n_1047) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_927), .A2(n_800), .B1(n_808), .B2(n_895), .C(n_814), .Y(n_1048) );
OAI221xp5_ASAP7_75t_SL g1049 ( .A1(n_924), .A2(n_880), .B1(n_907), .B2(n_889), .C(n_885), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_924), .A2(n_907), .B1(n_889), .B2(n_885), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1030), .Y(n_1051) );
OAI21xp5_ASAP7_75t_SL g1052 ( .A1(n_969), .A2(n_838), .B(n_859), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_954), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_911), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_925), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_973), .Y(n_1056) );
AOI31xp33_ASAP7_75t_L g1057 ( .A1(n_1004), .A2(n_825), .A3(n_838), .B(n_852), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_1035), .B(n_899), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_976), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_994), .B(n_798), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_973), .Y(n_1061) );
NOR2xp33_ASAP7_75t_R g1062 ( .A(n_982), .B(n_898), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1063 ( .A(n_938), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_948), .B(n_799), .Y(n_1064) );
AND4x1_ASAP7_75t_L g1065 ( .A(n_1002), .B(n_898), .C(n_153), .D(n_155), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_1001), .B(n_906), .C(n_891), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_991), .A2(n_825), .B1(n_891), .B2(n_864), .Y(n_1067) );
OAI321xp33_ASAP7_75t_L g1068 ( .A1(n_956), .A2(n_969), .A3(n_975), .B1(n_1015), .B2(n_999), .C(n_989), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_958), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_1035), .B(n_891), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_913), .Y(n_1071) );
AOI211xp5_ASAP7_75t_L g1072 ( .A1(n_979), .A2(n_891), .B(n_864), .C(n_865), .Y(n_1072) );
NAND4xp25_ASAP7_75t_L g1073 ( .A(n_997), .B(n_864), .C(n_865), .D(n_157), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_978), .B(n_864), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_910), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_914), .B(n_151), .Y(n_1076) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_1016), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_937), .B(n_156), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_985), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1006), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_991), .A2(n_158), .B1(n_159), .B2(n_161), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_958), .Y(n_1082) );
OAI31xp33_ASAP7_75t_SL g1083 ( .A1(n_1013), .A2(n_162), .A3(n_164), .B(n_165), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_1029), .A2(n_166), .B1(n_168), .B2(n_171), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_973), .Y(n_1085) );
INVx2_ASAP7_75t_L g1086 ( .A(n_945), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_965), .Y(n_1087) );
AOI22xp33_ASAP7_75t_SL g1088 ( .A1(n_1013), .A2(n_172), .B1(n_174), .B2(n_176), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_957), .B(n_177), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_945), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1003), .B(n_1023), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_944), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_956), .A2(n_186), .B1(n_188), .B2(n_189), .C(n_190), .Y(n_1093) );
AO21x2_ASAP7_75t_L g1094 ( .A1(n_1036), .A2(n_194), .B(n_197), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_918), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_962), .B(n_199), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_909), .A2(n_200), .B1(n_202), .B2(n_207), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_918), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_930), .A2(n_217), .B1(n_226), .B2(n_227), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_992), .B(n_229), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1005), .B(n_230), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_952), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1012), .B(n_233), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_909), .A2(n_234), .B1(n_236), .B2(n_237), .Y(n_1104) );
OA21x2_ASAP7_75t_L g1105 ( .A1(n_934), .A2(n_238), .B(n_239), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_1003), .B(n_240), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1019), .B(n_241), .Y(n_1107) );
AOI31xp33_ASAP7_75t_L g1108 ( .A1(n_1004), .A2(n_243), .A3(n_244), .B(n_245), .Y(n_1108) );
AOI211xp5_ASAP7_75t_L g1109 ( .A1(n_999), .A2(n_246), .B(n_248), .C(n_249), .Y(n_1109) );
NAND4xp25_ASAP7_75t_SL g1110 ( .A(n_981), .B(n_250), .C(n_251), .D(n_253), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_984), .A2(n_254), .B1(n_255), .B2(n_260), .C(n_262), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_995), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_960), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1023), .B(n_263), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_915), .B(n_264), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_974), .Y(n_1116) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_940), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_973), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_972), .A2(n_265), .B1(n_266), .B2(n_267), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_912), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_949), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1041), .Y(n_1122) );
NAND2xp33_ASAP7_75t_R g1123 ( .A(n_1034), .B(n_268), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_998), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_1020), .A2(n_269), .B1(n_270), .B2(n_272), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_993), .A2(n_273), .B1(n_277), .B2(n_278), .Y(n_1126) );
AO21x2_ASAP7_75t_L g1127 ( .A1(n_1036), .A2(n_280), .B(n_284), .Y(n_1127) );
NOR2xp33_ASAP7_75t_R g1128 ( .A(n_1032), .B(n_285), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_914), .B(n_286), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1018), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_964), .B(n_287), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_964), .B(n_288), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_966), .B(n_290), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_942), .A2(n_291), .B1(n_293), .B2(n_294), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1039), .Y(n_1135) );
AO21x2_ASAP7_75t_L g1136 ( .A1(n_1008), .A2(n_295), .B(n_297), .Y(n_1136) );
NOR2xp33_ASAP7_75t_R g1137 ( .A(n_916), .B(n_300), .Y(n_1137) );
NAND2xp33_ASAP7_75t_SL g1138 ( .A(n_1033), .B(n_939), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_921), .A2(n_928), .B1(n_1000), .B2(n_931), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1007), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_987), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_917), .Y(n_1142) );
INVx2_ASAP7_75t_L g1143 ( .A(n_966), .Y(n_1143) );
OAI21xp5_ASAP7_75t_L g1144 ( .A1(n_972), .A2(n_963), .B(n_971), .Y(n_1144) );
OAI21x1_ASAP7_75t_L g1145 ( .A1(n_986), .A2(n_935), .B(n_943), .Y(n_1145) );
NAND3xp33_ASAP7_75t_L g1146 ( .A(n_1014), .B(n_983), .C(n_996), .Y(n_1146) );
INVxp67_ASAP7_75t_L g1147 ( .A(n_1011), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_1139), .A2(n_1014), .B1(n_1009), .B2(n_988), .Y(n_1148) );
NOR3xp33_ASAP7_75t_L g1149 ( .A(n_1147), .B(n_959), .C(n_950), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1054), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1074), .B(n_1009), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_1146), .A2(n_1135), .B(n_1025), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1055), .Y(n_1153) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_1138), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1074), .Y(n_1155) );
INVx3_ASAP7_75t_L g1156 ( .A(n_1070), .Y(n_1156) );
INVx4_ASAP7_75t_L g1157 ( .A(n_1046), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1075), .Y(n_1158) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_1062), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1160 ( .A1(n_1141), .A2(n_950), .B1(n_1022), .B2(n_1015), .C(n_980), .Y(n_1160) );
INVx3_ASAP7_75t_L g1161 ( .A(n_1070), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1063), .B(n_929), .Y(n_1162) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1069), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1120), .B(n_1024), .Y(n_1164) );
AOI21xp33_ASAP7_75t_SL g1165 ( .A1(n_1108), .A2(n_990), .B(n_1021), .Y(n_1165) );
OAI21xp5_ASAP7_75t_L g1166 ( .A1(n_1135), .A2(n_988), .B(n_977), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1079), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1112), .B(n_959), .Y(n_1168) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1070), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1080), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1122), .Y(n_1171) );
NAND4xp25_ASAP7_75t_L g1172 ( .A(n_1060), .B(n_1017), .C(n_936), .D(n_970), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1056), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1056), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1042), .B(n_951), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1061), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1069), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1113), .B(n_919), .Y(n_1178) );
OAI21xp5_ASAP7_75t_SL g1179 ( .A1(n_1057), .A2(n_1033), .B(n_923), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1142), .B(n_1021), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1071), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1117), .B(n_951), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1047), .B(n_1051), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1087), .B(n_1021), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1053), .B(n_970), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1047), .B(n_953), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_1138), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_1110), .A2(n_961), .B1(n_932), .B2(n_936), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1051), .B(n_947), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1061), .B(n_946), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1059), .B(n_920), .Y(n_1191) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_1077), .Y(n_1192) );
OAI33xp33_ASAP7_75t_L g1193 ( .A1(n_1130), .A2(n_1028), .A3(n_1031), .B1(n_1026), .B2(n_951), .B3(n_1038), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1082), .Y(n_1194) );
AOI311xp33_ASAP7_75t_L g1195 ( .A1(n_1140), .A2(n_1028), .A3(n_986), .B(n_1037), .C(n_922), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1085), .B(n_955), .Y(n_1196) );
AOI31xp33_ASAP7_75t_L g1197 ( .A1(n_1123), .A2(n_941), .A3(n_926), .B(n_933), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1085), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1116), .B(n_941), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1118), .B(n_926), .Y(n_1200) );
BUFx2_ASAP7_75t_L g1201 ( .A(n_1117), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1118), .B(n_933), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1082), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1086), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1129), .Y(n_1205) );
BUFx3_ASAP7_75t_L g1206 ( .A(n_1046), .Y(n_1206) );
INVx4_ASAP7_75t_L g1207 ( .A(n_1076), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1121), .B(n_1040), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1121), .B(n_967), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1210 ( .A(n_1143), .Y(n_1210) );
NAND2x1p5_ASAP7_75t_L g1211 ( .A(n_1129), .B(n_967), .Y(n_1211) );
NAND2x1p5_ASAP7_75t_L g1212 ( .A(n_1133), .B(n_1106), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1042), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1045), .B(n_1095), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1045), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1143), .B(n_1102), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1064), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1091), .B(n_1052), .Y(n_1218) );
AOI22xp33_ASAP7_75t_SL g1219 ( .A1(n_1128), .A2(n_1131), .B1(n_1132), .B2(n_1137), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1091), .B(n_1132), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1133), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1102), .B(n_1086), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1131), .B(n_1043), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1072), .B(n_1083), .C(n_1065), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1106), .Y(n_1225) );
OAI33xp33_ASAP7_75t_L g1226 ( .A1(n_1073), .A2(n_1126), .A3(n_1050), .B1(n_1119), .B2(n_1098), .B3(n_1084), .Y(n_1226) );
INVx1_ASAP7_75t_SL g1227 ( .A(n_1076), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1090), .B(n_1107), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_1068), .A2(n_1093), .B1(n_1044), .B2(n_1144), .C(n_1067), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1090), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1124), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1107), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1170), .Y(n_1233) );
NOR2xp33_ASAP7_75t_R g1234 ( .A(n_1207), .B(n_1076), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1163), .Y(n_1235) );
AND3x1_ASAP7_75t_L g1236 ( .A(n_1185), .B(n_1109), .C(n_1111), .Y(n_1236) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1181), .B(n_1058), .Y(n_1237) );
NAND3xp33_ASAP7_75t_L g1238 ( .A(n_1149), .B(n_1088), .C(n_1104), .Y(n_1238) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_1182), .B(n_1145), .Y(n_1239) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1163), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1150), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1217), .B(n_1158), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1192), .B(n_1215), .Y(n_1243) );
CKINVDCx16_ASAP7_75t_R g1244 ( .A(n_1159), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1171), .B(n_1058), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1153), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1167), .Y(n_1247) );
NAND4xp25_ASAP7_75t_L g1248 ( .A(n_1219), .B(n_1097), .C(n_1099), .D(n_1081), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1155), .B(n_1145), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1213), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1172), .B(n_1115), .Y(n_1251) );
NAND2xp33_ASAP7_75t_R g1252 ( .A(n_1154), .B(n_1105), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1213), .Y(n_1253) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1229), .B(n_1066), .C(n_1048), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1216), .B(n_1058), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1214), .Y(n_1256) );
INVx4_ASAP7_75t_L g1257 ( .A(n_1207), .Y(n_1257) );
OR2x4_ASAP7_75t_L g1258 ( .A(n_1197), .B(n_1127), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1214), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1155), .Y(n_1260) );
OR2x6_ASAP7_75t_L g1261 ( .A(n_1207), .B(n_1114), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1200), .B(n_1103), .Y(n_1262) );
NOR2xp33_ASAP7_75t_R g1263 ( .A(n_1159), .B(n_1114), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1223), .B(n_1101), .Y(n_1264) );
INVx1_ASAP7_75t_SL g1265 ( .A(n_1184), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1162), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1173), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1173), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1164), .B(n_1101), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g1270 ( .A(n_1230), .Y(n_1270) );
NAND2x1_ASAP7_75t_L g1271 ( .A(n_1154), .B(n_1105), .Y(n_1271) );
OAI221xp5_ASAP7_75t_L g1272 ( .A1(n_1152), .A2(n_1134), .B1(n_1049), .B2(n_1092), .C(n_1125), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1200), .B(n_1078), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1228), .B(n_1105), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1151), .B(n_1078), .Y(n_1275) );
NOR3xp33_ASAP7_75t_SL g1276 ( .A(n_1179), .B(n_1094), .C(n_1127), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1174), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1151), .B(n_1089), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1218), .B(n_1089), .Y(n_1279) );
INVxp67_ASAP7_75t_L g1280 ( .A(n_1180), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1174), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1228), .B(n_1094), .Y(n_1282) );
INVx1_ASAP7_75t_SL g1283 ( .A(n_1206), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_1182), .B(n_1124), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1176), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1176), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1220), .B(n_1096), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1198), .Y(n_1288) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_1230), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1232), .B(n_1096), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_1157), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1177), .Y(n_1292) );
INVx2_ASAP7_75t_SL g1293 ( .A(n_1157), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1191), .B(n_1100), .Y(n_1294) );
NAND4xp25_ASAP7_75t_L g1295 ( .A(n_1224), .B(n_1100), .C(n_1094), .D(n_1127), .Y(n_1295) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1165), .B(n_1136), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1267), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1268), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1266), .B(n_1221), .Y(n_1299) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_1233), .A2(n_1148), .B1(n_1178), .B2(n_1168), .C(n_1201), .Y(n_1300) );
NAND3xp33_ASAP7_75t_L g1301 ( .A(n_1276), .B(n_1195), .C(n_1188), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1277), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_1248), .A2(n_1226), .B1(n_1187), .B2(n_1201), .Y(n_1303) );
AOI211xp5_ASAP7_75t_L g1304 ( .A1(n_1296), .A2(n_1187), .B(n_1182), .C(n_1227), .Y(n_1304) );
OAI31xp33_ASAP7_75t_L g1305 ( .A1(n_1251), .A2(n_1212), .A3(n_1205), .B(n_1206), .Y(n_1305) );
INVxp67_ASAP7_75t_L g1306 ( .A(n_1291), .Y(n_1306) );
OAI21xp5_ASAP7_75t_L g1307 ( .A1(n_1254), .A2(n_1166), .B(n_1160), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1242), .B(n_1222), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1260), .B(n_1222), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1249), .B(n_1202), .Y(n_1310) );
OAI21xp33_ASAP7_75t_L g1311 ( .A1(n_1276), .A2(n_1198), .B(n_1190), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1281), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_1251), .A2(n_1199), .B1(n_1193), .B2(n_1225), .C(n_1190), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1285), .Y(n_1314) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1244), .B(n_1157), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1256), .B(n_1202), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1280), .B(n_1175), .Y(n_1317) );
AOI322xp5_ASAP7_75t_L g1318 ( .A1(n_1296), .A2(n_1196), .A3(n_1209), .B1(n_1208), .B2(n_1183), .C1(n_1210), .C2(n_1204), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1249), .B(n_1196), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1286), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1282), .B(n_1183), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_1261), .A2(n_1212), .B1(n_1211), .B2(n_1175), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1259), .B(n_1209), .Y(n_1323) );
NOR2x1_ASAP7_75t_L g1324 ( .A(n_1257), .B(n_1156), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1241), .B(n_1210), .Y(n_1325) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_1261), .A2(n_1212), .B1(n_1211), .B2(n_1161), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1282), .B(n_1204), .Y(n_1327) );
AOI21xp5_ASAP7_75t_L g1328 ( .A1(n_1258), .A2(n_1211), .B(n_1208), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1288), .Y(n_1329) );
INVx1_ASAP7_75t_SL g1330 ( .A(n_1283), .Y(n_1330) );
AOI21xp5_ASAP7_75t_L g1331 ( .A1(n_1258), .A2(n_1136), .B(n_1203), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1274), .B(n_1203), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1274), .B(n_1177), .Y(n_1333) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1235), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1250), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1253), .Y(n_1336) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1235), .Y(n_1337) );
A2O1A1Ixp33_ASAP7_75t_L g1338 ( .A1(n_1291), .A2(n_1156), .B(n_1161), .C(n_1169), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_1261), .A2(n_1156), .B1(n_1161), .B2(n_1169), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_1279), .A2(n_1169), .B1(n_1186), .B2(n_1189), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1255), .B(n_1194), .Y(n_1341) );
OAI21xp5_ASAP7_75t_SL g1342 ( .A1(n_1303), .A2(n_1295), .B(n_1293), .Y(n_1342) );
NAND2xp33_ASAP7_75t_R g1343 ( .A(n_1315), .B(n_1234), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1297), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1310), .B(n_1239), .Y(n_1345) );
OAI32xp33_ASAP7_75t_L g1346 ( .A1(n_1330), .A2(n_1306), .A3(n_1257), .B1(n_1301), .B2(n_1265), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1310), .B(n_1243), .Y(n_1347) );
INVx1_ASAP7_75t_SL g1348 ( .A(n_1341), .Y(n_1348) );
INVxp33_ASAP7_75t_SL g1349 ( .A(n_1322), .Y(n_1349) );
NAND2xp33_ASAP7_75t_SL g1350 ( .A(n_1340), .B(n_1234), .Y(n_1350) );
INVx2_ASAP7_75t_SL g1351 ( .A(n_1324), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1319), .B(n_1247), .Y(n_1352) );
INVxp33_ASAP7_75t_L g1353 ( .A(n_1317), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1297), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1298), .Y(n_1355) );
NOR3xp33_ASAP7_75t_SL g1356 ( .A(n_1307), .B(n_1272), .C(n_1238), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1298), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1302), .Y(n_1358) );
CKINVDCx20_ASAP7_75t_R g1359 ( .A(n_1308), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1319), .B(n_1239), .Y(n_1360) );
HB1xp67_ASAP7_75t_L g1361 ( .A(n_1341), .Y(n_1361) );
NAND2xp33_ASAP7_75t_SL g1362 ( .A(n_1339), .B(n_1263), .Y(n_1362) );
NOR3xp33_ASAP7_75t_SL g1363 ( .A(n_1300), .B(n_1252), .C(n_1294), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1302), .Y(n_1364) );
NAND2x1_ASAP7_75t_L g1365 ( .A(n_1328), .B(n_1257), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1313), .B(n_1246), .C(n_1236), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1316), .B(n_1289), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1321), .B(n_1289), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1312), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1312), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1314), .Y(n_1371) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1334), .Y(n_1372) );
AOI322xp5_ASAP7_75t_L g1373 ( .A1(n_1362), .A2(n_1311), .A3(n_1326), .B1(n_1299), .B2(n_1321), .C1(n_1293), .C2(n_1323), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1366), .Y(n_1374) );
AOI211xp5_ASAP7_75t_L g1375 ( .A1(n_1346), .A2(n_1305), .B(n_1304), .C(n_1263), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_1349), .A2(n_1252), .B1(n_1269), .B2(n_1325), .Y(n_1376) );
OAI32xp33_ASAP7_75t_L g1377 ( .A1(n_1349), .A2(n_1237), .A3(n_1309), .B1(n_1270), .B2(n_1245), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1367), .B(n_1318), .Y(n_1378) );
NOR2x1_ASAP7_75t_L g1379 ( .A(n_1365), .B(n_1338), .Y(n_1379) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1372), .Y(n_1380) );
OAI211xp5_ASAP7_75t_L g1381 ( .A1(n_1356), .A2(n_1331), .B(n_1264), .C(n_1290), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1345), .B(n_1327), .Y(n_1382) );
NAND4xp25_ASAP7_75t_SL g1383 ( .A(n_1359), .B(n_1278), .C(n_1275), .D(n_1273), .Y(n_1383) );
NAND2xp5_ASAP7_75t_SL g1384 ( .A(n_1362), .B(n_1270), .Y(n_1384) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1372), .Y(n_1385) );
AOI211xp5_ASAP7_75t_L g1386 ( .A1(n_1346), .A2(n_1239), .B(n_1336), .C(n_1335), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1370), .Y(n_1387) );
BUFx2_ASAP7_75t_L g1388 ( .A(n_1351), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1370), .Y(n_1389) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1361), .Y(n_1390) );
XNOR2xp5_ASAP7_75t_L g1391 ( .A(n_1359), .B(n_1287), .Y(n_1391) );
NAND2xp5_ASAP7_75t_SL g1392 ( .A(n_1350), .B(n_1284), .Y(n_1392) );
NAND3x1_ASAP7_75t_SL g1393 ( .A(n_1379), .B(n_1350), .C(n_1365), .Y(n_1393) );
OAI21xp5_ASAP7_75t_L g1394 ( .A1(n_1374), .A2(n_1342), .B(n_1363), .Y(n_1394) );
NOR3xp33_ASAP7_75t_L g1395 ( .A(n_1381), .B(n_1384), .C(n_1392), .Y(n_1395) );
INVx2_ASAP7_75t_SL g1396 ( .A(n_1388), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1387), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1382), .B(n_1345), .Y(n_1398) );
OAI221xp5_ASAP7_75t_L g1399 ( .A1(n_1373), .A2(n_1351), .B1(n_1343), .B2(n_1353), .C(n_1348), .Y(n_1399) );
NOR2xp33_ASAP7_75t_R g1400 ( .A(n_1383), .B(n_1347), .Y(n_1400) );
A2O1A1Ixp33_ASAP7_75t_L g1401 ( .A1(n_1373), .A2(n_1360), .B(n_1368), .C(n_1352), .Y(n_1401) );
AOI321xp33_ASAP7_75t_L g1402 ( .A1(n_1375), .A2(n_1360), .A3(n_1369), .B1(n_1364), .B2(n_1371), .C(n_1358), .Y(n_1402) );
XNOR2xp5_ASAP7_75t_L g1403 ( .A(n_1391), .B(n_1262), .Y(n_1403) );
OAI22x1_ASAP7_75t_L g1404 ( .A1(n_1391), .A2(n_1357), .B1(n_1355), .B2(n_1354), .Y(n_1404) );
INVx2_ASAP7_75t_L g1405 ( .A(n_1390), .Y(n_1405) );
AO22x2_ASAP7_75t_L g1406 ( .A1(n_1378), .A2(n_1344), .B1(n_1314), .B2(n_1320), .Y(n_1406) );
OAI222xp33_ASAP7_75t_L g1407 ( .A1(n_1379), .A2(n_1336), .B1(n_1335), .B2(n_1320), .C1(n_1329), .C2(n_1327), .Y(n_1407) );
OAI211xp5_ASAP7_75t_L g1408 ( .A1(n_1386), .A2(n_1329), .B(n_1271), .C(n_1332), .Y(n_1408) );
OA22x2_ASAP7_75t_L g1409 ( .A1(n_1388), .A2(n_1333), .B1(n_1332), .B2(n_1284), .Y(n_1409) );
NOR3xp33_ASAP7_75t_L g1410 ( .A(n_1376), .B(n_1337), .C(n_1334), .Y(n_1410) );
AOI211xp5_ASAP7_75t_L g1411 ( .A1(n_1377), .A2(n_1284), .B(n_1186), .C(n_1189), .Y(n_1411) );
XOR2xp5_ASAP7_75t_L g1412 ( .A(n_1382), .B(n_1240), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_1389), .A2(n_1292), .B1(n_1136), .B2(n_1194), .Y(n_1413) );
NAND4xp75_ASAP7_75t_L g1414 ( .A(n_1387), .B(n_1231), .C(n_1292), .D(n_1389), .Y(n_1414) );
INVx1_ASAP7_75t_SL g1415 ( .A(n_1396), .Y(n_1415) );
NOR2x1p5_ASAP7_75t_L g1416 ( .A(n_1393), .B(n_1414), .Y(n_1416) );
OAI221xp5_ASAP7_75t_R g1417 ( .A1(n_1403), .A2(n_1395), .B1(n_1399), .B2(n_1410), .C(n_1412), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1397), .Y(n_1418) );
NAND3xp33_ASAP7_75t_SL g1419 ( .A(n_1394), .B(n_1399), .C(n_1402), .Y(n_1419) );
NOR2xp67_ASAP7_75t_L g1420 ( .A(n_1408), .B(n_1404), .Y(n_1420) );
AOI22xp33_ASAP7_75t_SL g1421 ( .A1(n_1417), .A2(n_1394), .B1(n_1406), .B2(n_1400), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1415), .B(n_1406), .Y(n_1422) );
XNOR2x1_ASAP7_75t_L g1423 ( .A(n_1416), .B(n_1409), .Y(n_1423) );
NAND4xp25_ASAP7_75t_L g1424 ( .A(n_1419), .B(n_1402), .C(n_1401), .D(n_1411), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1418), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1425), .Y(n_1426) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1422), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1423), .Y(n_1428) );
XNOR2xp5_ASAP7_75t_L g1429 ( .A(n_1421), .B(n_1420), .Y(n_1429) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1426), .Y(n_1430) );
INVxp67_ASAP7_75t_SL g1431 ( .A(n_1428), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_1429), .A2(n_1418), .B1(n_1424), .B2(n_1411), .Y(n_1432) );
AOI322xp5_ASAP7_75t_L g1433 ( .A1(n_1431), .A2(n_1427), .A3(n_1429), .B1(n_1405), .B2(n_1398), .C1(n_1413), .C2(n_1380), .Y(n_1433) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_1432), .A2(n_1427), .B1(n_1380), .B2(n_1385), .Y(n_1434) );
INVxp67_ASAP7_75t_L g1435 ( .A(n_1430), .Y(n_1435) );
AOI221xp5_ASAP7_75t_SL g1436 ( .A1(n_1435), .A2(n_1433), .B1(n_1434), .B2(n_1377), .C(n_1407), .Y(n_1436) );
endmodule