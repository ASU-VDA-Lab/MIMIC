module fake_jpeg_27994_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_27),
.B1(n_17),
.B2(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_65),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_21),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_24),
.C(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_74),
.Y(n_99)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_77),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_44),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_20),
.B1(n_22),
.B2(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_106),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_20),
.B(n_33),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_113),
.B(n_99),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_35),
.B1(n_63),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_109),
.B1(n_84),
.B2(n_82),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_20),
.A3(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_35),
.B1(n_38),
.B2(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_71),
.B1(n_78),
.B2(n_89),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_18),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_80),
.B1(n_72),
.B2(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_70),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_35),
.B1(n_51),
.B2(n_31),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_34),
.B(n_38),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_34),
.B(n_23),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_0),
.B(n_1),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_134),
.B1(n_139),
.B2(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_130),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_26),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_18),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_135),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_92),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_36),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_136),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_85),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_90),
.C(n_86),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_146),
.C(n_36),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_86),
.B1(n_83),
.B2(n_76),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_69),
.B1(n_34),
.B2(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_24),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_69),
.B1(n_16),
.B2(n_23),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_26),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_101),
.B(n_111),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_100),
.B(n_107),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_39),
.C(n_36),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_103),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_103),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_160),
.B(n_161),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_119),
.B(n_117),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_145),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_165),
.B(n_177),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_167),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_122),
.B(n_127),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_115),
.C(n_107),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_121),
.C(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_178),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_100),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_34),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_128),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_128),
.B1(n_145),
.B2(n_134),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_200),
.B1(n_202),
.B2(n_205),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_186),
.C(n_187),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_166),
.C(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_126),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_142),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_201),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_126),
.A3(n_147),
.B1(n_115),
.B2(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_120),
.B1(n_118),
.B2(n_102),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_206),
.B1(n_154),
.B2(n_178),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_207),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_120),
.B1(n_26),
.B2(n_23),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_34),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_16),
.B1(n_23),
.B2(n_26),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_24),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_26),
.B1(n_23),
.B2(n_16),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_151),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_34),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_229),
.Y(n_249)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_177),
.B1(n_161),
.B2(n_160),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_214),
.B1(n_222),
.B2(n_231),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_169),
.B(n_152),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_223),
.B(n_227),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_230),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_172),
.B1(n_179),
.B2(n_149),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_9),
.Y(n_252)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_162),
.C(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.C(n_199),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_159),
.C(n_156),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_156),
.B1(n_154),
.B2(n_176),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_31),
.B(n_11),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_186),
.B(n_31),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_9),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_185),
.B(n_184),
.C(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_203),
.B1(n_195),
.B2(n_182),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_29),
.B1(n_10),
.B2(n_15),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_236),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_221),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_227),
.B(n_209),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_201),
.B1(n_207),
.B2(n_2),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_250),
.B1(n_247),
.B2(n_213),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_29),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_41),
.C(n_39),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_41),
.C(n_39),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_0),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_41),
.C(n_39),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_252),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_215),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_216),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_257),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_211),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_233),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_223),
.C(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_227),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_0),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_237),
.B1(n_246),
.B2(n_241),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_269),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_254),
.A2(n_248),
.B(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_275),
.B1(n_279),
.B2(n_11),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_249),
.B1(n_233),
.B2(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_242),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_281),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_251),
.B1(n_253),
.B2(n_215),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_11),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_288),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_264),
.C(n_255),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_295),
.C(n_39),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_257),
.B1(n_269),
.B2(n_1),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_276),
.B(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_6),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_8),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_294),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_270),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_8),
.B(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_6),
.B(n_7),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_2),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_6),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_41),
.C(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_13),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_293),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_296),
.A2(n_286),
.B1(n_295),
.B2(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_300),
.B(n_14),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_305),
.B(n_306),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.B1(n_314),
.B2(n_310),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_307),
.C(n_13),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_13),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_41),
.Y(n_319)
);


endmodule