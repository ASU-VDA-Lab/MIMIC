module fake_jpeg_31510_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_34),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_54),
.B1(n_46),
.B2(n_50),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_50),
.C(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_16),
.B1(n_37),
.B2(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_39),
.B1(n_13),
.B2(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_3),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_12),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_8),
.C(n_9),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_27),
.C(n_26),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_103),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_105),
.B(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_24),
.C(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_94),
.B1(n_90),
.B2(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_112),
.B1(n_108),
.B2(n_106),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_114),
.B(n_104),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_103),
.C(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_115),
.B1(n_107),
.B2(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_113),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_120),
.Y(n_123)
);

OAI31xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_114),
.A3(n_99),
.B(n_116),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_99),
.C(n_9),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_18),
.B(n_20),
.Y(n_126)
);


endmodule