module fake_jpeg_4808_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_30),
.B(n_19),
.C(n_28),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_55),
.Y(n_82)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_56),
.B1(n_37),
.B2(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_17),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx2_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_50),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_69),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_40),
.B1(n_24),
.B2(n_23),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_23),
.B(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_38),
.B1(n_35),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_73),
.B1(n_50),
.B2(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_21),
.B1(n_38),
.B2(n_17),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_42),
.B1(n_79),
.B2(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_17),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_75),
.C(n_62),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_117),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2x1_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_72),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_98),
.B(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_84),
.B(n_66),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_63),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_72),
.C(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_46),
.B1(n_47),
.B2(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_84),
.A3(n_104),
.B1(n_94),
.B2(n_85),
.C1(n_98),
.C2(n_95),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_120),
.C(n_16),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_138),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_108),
.B(n_119),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_113),
.B1(n_123),
.B2(n_118),
.C(n_117),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_8),
.B(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_105),
.B1(n_121),
.B2(n_113),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_146),
.B1(n_138),
.B2(n_125),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_114),
.B1(n_123),
.B2(n_106),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_151),
.B(n_156),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_132),
.C(n_135),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_46),
.B1(n_90),
.B2(n_47),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_1),
.B(n_2),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_47),
.B1(n_89),
.B2(n_8),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_166),
.CI(n_148),
.CON(n_177),
.SN(n_177)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_140),
.C(n_136),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_167),
.C(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_164),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_130),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_149),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

XOR2x1_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_164),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_147),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_152),
.B1(n_129),
.B2(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_177),
.B(n_163),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_150),
.C(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_9),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_170),
.B1(n_160),
.B2(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_188),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_174),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_11),
.B1(n_9),
.B2(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_191),
.Y(n_198)
);

AOI31xp33_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_180),
.A3(n_178),
.B(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.C(n_2),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_185),
.C(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_4),
.C(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_189),
.C(n_6),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.C(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_5),
.C(n_6),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_202),
.Y(n_203)
);


endmodule