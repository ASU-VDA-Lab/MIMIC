module fake_aes_9194_n_1550 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1550);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1550;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1542;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVxp33_ASAP7_75t_SL g338 ( .A(n_323), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_194), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_267), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_12), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_219), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_74), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_310), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_57), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_193), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_116), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_190), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_264), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_166), .Y(n_350) );
INVxp33_ASAP7_75t_SL g351 ( .A(n_162), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_247), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_107), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_137), .Y(n_355) );
BUFx2_ASAP7_75t_SL g356 ( .A(n_55), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_86), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_152), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_97), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_318), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_76), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_204), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_201), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_39), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_246), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_53), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_135), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_31), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_257), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_82), .B(n_163), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_77), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_136), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_54), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_231), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_286), .Y(n_377) );
CKINVDCx14_ASAP7_75t_R g378 ( .A(n_141), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_93), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_28), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_75), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_183), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_203), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_108), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_131), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_303), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_0), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_87), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_146), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_66), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_270), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_79), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_202), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_125), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_112), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_327), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_199), .Y(n_397) );
CKINVDCx14_ASAP7_75t_R g398 ( .A(n_328), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_139), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_74), .Y(n_400) );
INVxp33_ASAP7_75t_L g401 ( .A(n_43), .Y(n_401) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_290), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_262), .Y(n_403) );
INVxp33_ASAP7_75t_SL g404 ( .A(n_189), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_43), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_59), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_69), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_113), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_311), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_331), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_226), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_20), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_20), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_276), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_12), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_248), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_288), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_8), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_106), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_260), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_317), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_238), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_15), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_79), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_245), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_313), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_161), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_195), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_232), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_147), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_225), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_29), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_191), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_237), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_93), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_322), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_165), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_261), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_334), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_76), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_312), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_263), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_298), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_206), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_36), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_205), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_182), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_89), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_18), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_96), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_1), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_159), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_5), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_34), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_30), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_239), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_21), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_250), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_95), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_251), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_181), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_255), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_266), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_207), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_269), .Y(n_465) );
INVxp33_ASAP7_75t_SL g466 ( .A(n_240), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_31), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_68), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_34), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_39), .Y(n_470) );
INVxp33_ASAP7_75t_SL g471 ( .A(n_138), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_96), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_58), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_41), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_71), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_28), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_287), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_271), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_89), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_126), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_25), .Y(n_481) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_293), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_301), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_198), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_27), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_101), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_112), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_98), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_122), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_282), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_309), .Y(n_491) );
INVxp33_ASAP7_75t_SL g492 ( .A(n_111), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_95), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_35), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_117), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_324), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_111), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_325), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_285), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_37), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_299), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_227), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_273), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_321), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_346), .B(n_0), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_383), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_383), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_345), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_346), .B(n_384), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_444), .B(n_1), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_396), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_376), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_345), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_385), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_385), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_444), .B(n_2), .Y(n_517) );
AND3x2_ASAP7_75t_L g518 ( .A(n_475), .B(n_2), .C(n_3), .Y(n_518) );
NAND2xp33_ASAP7_75t_L g519 ( .A(n_412), .B(n_124), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_386), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_386), .Y(n_521) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_396), .A2(n_128), .B(n_127), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_376), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_376), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_389), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_401), .B(n_3), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_379), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_389), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_376), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_376), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_419), .B(n_4), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_373), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_384), .B(n_4), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_399), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_388), .B(n_5), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_399), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_391), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_391), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_436), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_365), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_410), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_379), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_388), .B(n_6), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_508), .B(n_344), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_508), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_508), .B(n_431), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_527), .B(n_425), .Y(n_547) );
NAND3x1_ASAP7_75t_L g548 ( .A(n_533), .B(n_392), .C(n_390), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_527), .B(n_439), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_513), .B(n_378), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_511), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_527), .B(n_410), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_341), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_513), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_511), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_511), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_532), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_514), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_514), .B(n_398), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_523), .Y(n_567) );
INVx4_ASAP7_75t_L g568 ( .A(n_510), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_510), .B(n_452), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_523), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_533), .B(n_468), .C(n_423), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_506), .B(n_452), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_509), .B(n_461), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_511), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_533), .B(n_356), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_526), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_523), .Y(n_580) );
INVx5_ASAP7_75t_L g581 ( .A(n_523), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_509), .B(n_491), .Y(n_582) );
AND2x6_ASAP7_75t_L g583 ( .A(n_510), .B(n_517), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_534), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_534), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_534), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_542), .B(n_442), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_510), .B(n_424), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_524), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_568), .B(n_517), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_574), .B(n_509), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_574), .B(n_542), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_582), .B(n_526), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_579), .Y(n_597) );
AND2x6_ASAP7_75t_L g598 ( .A(n_557), .B(n_517), .Y(n_598) );
INVx4_ASAP7_75t_L g599 ( .A(n_583), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_569), .A2(n_522), .B(n_517), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
INVx5_ASAP7_75t_L g603 ( .A(n_583), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
OR2x6_ASAP7_75t_L g605 ( .A(n_556), .B(n_531), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_571), .Y(n_608) );
BUFx4f_ASAP7_75t_L g609 ( .A(n_577), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_552), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_582), .B(n_526), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_583), .A2(n_507), .B1(n_515), .B2(n_506), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_545), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_577), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_555), .A2(n_374), .B1(n_420), .B2(n_349), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_545), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_568), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_583), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_507), .B1(n_515), .B2(n_506), .Y(n_620) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_557), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_568), .B(n_517), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_547), .B(n_531), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_556), .B(n_531), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_577), .Y(n_626) );
INVx4_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_557), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_577), .Y(n_629) );
INVx5_ASAP7_75t_L g630 ( .A(n_583), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_577), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_568), .B(n_507), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_552), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_556), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_547), .B(n_531), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_577), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_589), .Y(n_637) );
BUFx3_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_549), .B(n_515), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_544), .A2(n_505), .B1(n_492), .B2(n_374), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_589), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_589), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_549), .B(n_505), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_588), .B(n_516), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_554), .B(n_516), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_562), .Y(n_648) );
OR2x6_ASAP7_75t_L g649 ( .A(n_555), .B(n_356), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_583), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_544), .A2(n_492), .B1(n_420), .B2(n_434), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_551), .Y(n_652) );
BUFx3_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_551), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_564), .B(n_535), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_583), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_588), .B(n_516), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_558), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_555), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_588), .B(n_520), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_544), .A2(n_434), .B1(n_462), .B2(n_349), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_550), .B(n_520), .Y(n_665) );
BUFx4f_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_559), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_546), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_560), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_568), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_546), .A2(n_572), .B1(n_550), .B2(n_565), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_546), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_552), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_560), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_554), .B(n_520), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_561), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_562), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_591), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_591), .B(n_521), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_561), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_591), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_576), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_589), .Y(n_683) );
NOR2x1p5_ASAP7_75t_L g684 ( .A(n_565), .B(n_341), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_565), .B(n_521), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_589), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_576), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_686), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_683), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_594), .B(n_572), .Y(n_690) );
INVx5_ASAP7_75t_L g691 ( .A(n_650), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_660), .A2(n_462), .B1(n_548), .B2(n_589), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_647), .B(n_591), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_671), .B(n_569), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_683), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_686), .Y(n_696) );
BUFx3_ASAP7_75t_L g697 ( .A(n_613), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_683), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_596), .B(n_591), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_647), .B(n_548), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_597), .B(n_518), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_602), .A2(n_548), .B1(n_343), .B2(n_407), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_616), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_683), .Y(n_704) );
AND2x4_ASAP7_75t_SL g705 ( .A(n_605), .B(n_532), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_605), .B(n_373), .Y(n_706) );
BUFx3_ASAP7_75t_L g707 ( .A(n_668), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_686), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_617), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_600), .B(n_518), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_604), .B(n_535), .Y(n_711) );
NAND2x1_ASAP7_75t_L g712 ( .A(n_598), .B(n_578), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_617), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_609), .A2(n_573), .B1(n_525), .B2(n_528), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_655), .Y(n_715) );
INVx5_ASAP7_75t_L g716 ( .A(n_650), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_617), .Y(n_717) );
NAND2x1_ASAP7_75t_SL g718 ( .A(n_662), .B(n_405), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_637), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_675), .A2(n_573), .B(n_525), .C(n_528), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_675), .B(n_578), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_668), .Y(n_722) );
NAND2xp5_ASAP7_75t_R g723 ( .A(n_651), .B(n_405), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_650), .Y(n_724) );
INVx5_ASAP7_75t_L g725 ( .A(n_650), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_637), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_634), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_607), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_601), .A2(n_522), .B(n_519), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_605), .B(n_448), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_599), .B(n_584), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_643), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_624), .B(n_448), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_609), .A2(n_525), .B1(n_528), .B2(n_521), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_612), .A2(n_538), .B1(n_537), .B2(n_584), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_643), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_603), .Y(n_737) );
OR2x6_ASAP7_75t_L g738 ( .A(n_615), .B(n_535), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_644), .Y(n_739) );
BUFx2_ASAP7_75t_L g740 ( .A(n_634), .Y(n_740) );
BUFx4_ASAP7_75t_SL g741 ( .A(n_624), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_644), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_611), .B(n_587), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_603), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_610), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_612), .A2(n_538), .B1(n_537), .B2(n_587), .Y(n_746) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_603), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_606), .A2(n_543), .B1(n_540), .B2(n_538), .C(n_537), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_624), .Y(n_749) );
OR2x2_ASAP7_75t_SL g750 ( .A(n_648), .B(n_479), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_649), .A2(n_543), .B1(n_485), .B2(n_479), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_648), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_672), .A2(n_343), .B1(n_407), .B2(n_362), .Y(n_753) );
INVxp67_ASAP7_75t_L g754 ( .A(n_649), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_608), .B(n_543), .Y(n_755) );
BUFx2_ASAP7_75t_L g756 ( .A(n_649), .Y(n_756) );
NOR2xp33_ASAP7_75t_R g757 ( .A(n_677), .B(n_485), .Y(n_757) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_603), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_639), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_630), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_666), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_630), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g763 ( .A1(n_645), .A2(n_522), .B(n_536), .C(n_534), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_666), .B(n_362), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_630), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_684), .B(n_380), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_642), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_607), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_641), .B(n_454), .Y(n_769) );
BUFx2_ASAP7_75t_L g770 ( .A(n_677), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_610), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_619), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_598), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_595), .B(n_338), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_619), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_645), .Y(n_776) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_630), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_607), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_646), .B(n_454), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_658), .B(n_455), .Y(n_780) );
BUFx10_ASAP7_75t_L g781 ( .A(n_614), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_607), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_685), .B(n_400), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_633), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_618), .Y(n_785) );
CKINVDCx8_ASAP7_75t_R g786 ( .A(n_598), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_661), .B(n_347), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_625), .B(n_354), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_652), .Y(n_789) );
INVx4_ASAP7_75t_L g790 ( .A(n_598), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_620), .A2(n_536), .B1(n_541), .B2(n_534), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_598), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_593), .A2(n_522), .B(n_519), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_626), .B(n_357), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_618), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_621), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_633), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_623), .Y(n_798) );
INVx4_ASAP7_75t_L g799 ( .A(n_621), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_654), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_621), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_629), .A2(n_473), .B1(n_474), .B2(n_455), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_631), .A2(n_474), .B1(n_476), .B2(n_473), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_656), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_659), .Y(n_805) );
BUFx12f_ASAP7_75t_L g806 ( .A(n_599), .Y(n_806) );
OR2x6_ASAP7_75t_L g807 ( .A(n_638), .B(n_390), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_L g808 ( .A1(n_665), .A2(n_540), .B(n_489), .C(n_392), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_599), .B(n_424), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_636), .A2(n_488), .B1(n_476), .B2(n_351), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_638), .Y(n_811) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_653), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_627), .A2(n_541), .B1(n_536), .B2(n_351), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_627), .A2(n_541), .B1(n_536), .B2(n_404), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_621), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_628), .Y(n_816) );
BUFx12f_ASAP7_75t_L g817 ( .A(n_627), .Y(n_817) );
INVx3_ASAP7_75t_L g818 ( .A(n_628), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_663), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_620), .A2(n_640), .B1(n_657), .B2(n_653), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_664), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_635), .A2(n_488), .B1(n_404), .B2(n_466), .Y(n_822) );
INVx2_ASAP7_75t_SL g823 ( .A(n_657), .Y(n_823) );
OR2x6_ASAP7_75t_L g824 ( .A(n_593), .B(n_489), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_628), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_656), .Y(n_826) );
INVx2_ASAP7_75t_SL g827 ( .A(n_670), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_670), .B(n_338), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_667), .Y(n_829) );
NOR2x1_ASAP7_75t_L g830 ( .A(n_669), .B(n_497), .Y(n_830) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_628), .Y(n_831) );
BUFx2_ASAP7_75t_L g832 ( .A(n_687), .Y(n_832) );
AO31x2_ASAP7_75t_L g833 ( .A1(n_763), .A2(n_529), .A3(n_530), .B(n_512), .Y(n_833) );
AOI221x1_ASAP7_75t_L g834 ( .A1(n_763), .A2(n_540), .B1(n_350), .B2(n_352), .C(n_348), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_715), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_788), .Y(n_836) );
AO31x2_ASAP7_75t_L g837 ( .A1(n_729), .A2(n_529), .A3(n_530), .B(n_512), .Y(n_837) );
BUFx3_ASAP7_75t_L g838 ( .A(n_691), .Y(n_838) );
AND2x6_ASAP7_75t_L g839 ( .A(n_812), .B(n_673), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_776), .B(n_497), .Y(n_840) );
NOR2x1_ASAP7_75t_R g841 ( .A(n_752), .B(n_340), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_788), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_729), .A2(n_622), .B(n_679), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_SL g844 ( .A1(n_720), .A2(n_622), .B(n_353), .C(n_355), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_694), .A2(n_679), .B1(n_678), .B2(n_673), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_722), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_690), .A2(n_632), .B1(n_676), .B2(n_680), .C(n_674), .Y(n_847) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_705), .A2(n_471), .B1(n_466), .B2(n_368), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_694), .A2(n_681), .B1(n_678), .B2(n_682), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_789), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_706), .B(n_632), .Y(n_851) );
AO21x2_ASAP7_75t_L g852 ( .A1(n_793), .A2(n_529), .B(n_512), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_741), .Y(n_853) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_757), .A2(n_471), .B1(n_370), .B2(n_375), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_734), .A2(n_681), .B1(n_482), .B2(n_340), .Y(n_855) );
A2O1A1Ixp33_ASAP7_75t_L g856 ( .A1(n_699), .A2(n_541), .B(n_536), .C(n_365), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_745), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_798), .B(n_359), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_722), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_751), .A2(n_342), .B1(n_363), .B2(n_361), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_794), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_690), .A2(n_487), .B1(n_412), .B2(n_536), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_700), .A2(n_487), .B1(n_412), .B2(n_541), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_734), .A2(n_342), .B1(n_363), .B2(n_361), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_794), .Y(n_865) );
OAI211xp5_ASAP7_75t_L g866 ( .A1(n_718), .A2(n_381), .B(n_406), .C(n_395), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_824), .A2(n_377), .B1(n_421), .B2(n_364), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_771), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_738), .B(n_408), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_824), .A2(n_377), .B1(n_421), .B2(n_364), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_800), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_700), .A2(n_412), .B1(n_487), .B2(n_541), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_824), .A2(n_498), .B1(n_502), .B2(n_428), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_805), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_738), .A2(n_412), .B1(n_487), .B2(n_415), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_819), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_821), .Y(n_877) );
OAI222xp33_ASAP7_75t_L g878 ( .A1(n_751), .A2(n_500), .B1(n_481), .B2(n_486), .C1(n_472), .C2(n_432), .Y(n_878) );
INVx8_ASAP7_75t_L g879 ( .A(n_807), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_711), .B(n_413), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_829), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_772), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_714), .A2(n_498), .B1(n_502), .B2(n_428), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_759), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_786), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_767), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_738), .B(n_418), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_730), .B(n_440), .Y(n_888) );
INVx4_ASAP7_75t_L g889 ( .A(n_790), .Y(n_889) );
INVx4_ASAP7_75t_L g890 ( .A(n_790), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_711), .B(n_445), .Y(n_891) );
OAI22xp33_ASAP7_75t_L g892 ( .A1(n_692), .A2(n_435), .B1(n_457), .B2(n_387), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_775), .Y(n_893) );
AND2x6_ASAP7_75t_L g894 ( .A(n_812), .B(n_490), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_714), .A2(n_435), .B1(n_457), .B2(n_387), .Y(n_895) );
AND2x4_ASAP7_75t_L g896 ( .A(n_754), .B(n_449), .Y(n_896) );
OR2x6_ASAP7_75t_L g897 ( .A(n_741), .B(n_459), .Y(n_897) );
NAND2xp33_ASAP7_75t_L g898 ( .A(n_724), .B(n_436), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_784), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_807), .A2(n_456), .B1(n_496), .B2(n_402), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_797), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_755), .B(n_450), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_804), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_807), .A2(n_504), .B1(n_453), .B2(n_467), .Y(n_904) );
A2O1A1Ixp33_ASAP7_75t_L g905 ( .A1(n_699), .A2(n_470), .B(n_459), .C(n_469), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_826), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_755), .A2(n_487), .B1(n_493), .B2(n_451), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_697), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_820), .A2(n_495), .B1(n_494), .B2(n_470), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_820), .A2(n_458), .B1(n_358), .B2(n_360), .Y(n_910) );
AND2x4_ASAP7_75t_L g911 ( .A(n_754), .B(n_339), .Y(n_911) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_774), .A2(n_372), .B1(n_369), .B2(n_371), .C(n_367), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_783), .A2(n_382), .B1(n_393), .B2(n_366), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_831), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_703), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_832), .Y(n_916) );
AO21x2_ASAP7_75t_L g917 ( .A1(n_793), .A2(n_529), .B(n_512), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g918 ( .A1(n_757), .A2(n_397), .B1(n_443), .B2(n_414), .Y(n_918) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_749), .A2(n_397), .B1(n_443), .B2(n_414), .Y(n_919) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_779), .A2(n_480), .B1(n_446), .B2(n_403), .Y(n_920) );
INVx3_ASAP7_75t_L g921 ( .A(n_806), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_825), .Y(n_922) );
INVx2_ASAP7_75t_SL g923 ( .A(n_707), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_733), .B(n_6), .Y(n_924) );
OAI21x1_ASAP7_75t_L g925 ( .A1(n_809), .A2(n_830), .B(n_712), .Y(n_925) );
NOR2xp67_ASAP7_75t_L g926 ( .A(n_701), .B(n_7), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_727), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_779), .B(n_394), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_787), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_721), .A2(n_411), .B1(n_416), .B2(n_409), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_770), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_721), .A2(n_813), .B1(n_814), .B2(n_693), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_787), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_709), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_740), .B(n_7), .Y(n_935) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_724), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_783), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_764), .B(n_8), .Y(n_938) );
AND2x2_ASAP7_75t_SL g939 ( .A(n_756), .B(n_490), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_780), .B(n_417), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_761), .B(n_422), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_713), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_773), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_780), .B(n_426), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_693), .A2(n_566), .B(n_553), .Y(n_945) );
INVx2_ASAP7_75t_SL g946 ( .A(n_701), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_774), .B(n_427), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_748), .A2(n_430), .B1(n_433), .B2(n_429), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_831), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_769), .A2(n_480), .B1(n_446), .B2(n_437), .Y(n_950) );
BUFx2_ASAP7_75t_R g951 ( .A(n_792), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_766), .A2(n_465), .B1(n_438), .B2(n_447), .C(n_460), .Y(n_952) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_702), .A2(n_464), .B(n_477), .C(n_463), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_753), .B(n_9), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_822), .B(n_9), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_766), .A2(n_483), .B1(n_484), .B2(n_478), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_710), .B(n_499), .Y(n_957) );
BUFx12f_ASAP7_75t_L g958 ( .A(n_750), .Y(n_958) );
BUFx2_ASAP7_75t_L g959 ( .A(n_817), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_748), .B(n_503), .Y(n_960) );
A2O1A1Ixp33_ASAP7_75t_L g961 ( .A1(n_720), .A2(n_501), .B(n_530), .C(n_441), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_802), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_688), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_744), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_813), .A2(n_501), .B1(n_530), .B2(n_441), .Y(n_965) );
INVx2_ASAP7_75t_SL g966 ( .A(n_710), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_814), .A2(n_441), .B1(n_436), .B2(n_524), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_828), .A2(n_441), .B1(n_436), .B2(n_524), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_735), .A2(n_441), .B1(n_436), .B2(n_524), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_735), .B(n_10), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_746), .A2(n_13), .B1(n_10), .B2(n_11), .Y(n_971) );
OAI22x1_ASAP7_75t_L g972 ( .A1(n_723), .A2(n_14), .B1(n_11), .B2(n_13), .Y(n_972) );
INVx3_ASAP7_75t_L g973 ( .A(n_744), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_696), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_810), .B(n_14), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_803), .B(n_15), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_746), .A2(n_539), .B1(n_524), .B2(n_553), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_808), .A2(n_524), .B1(n_539), .B2(n_567), .C(n_580), .Y(n_978) );
OR2x6_ASAP7_75t_L g979 ( .A(n_795), .B(n_16), .Y(n_979) );
INVx2_ASAP7_75t_SL g980 ( .A(n_781), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_743), .A2(n_539), .B1(n_524), .B2(n_553), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_708), .Y(n_982) );
BUFx3_ASAP7_75t_L g983 ( .A(n_691), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_743), .A2(n_539), .B1(n_524), .B2(n_18), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_791), .Y(n_985) );
NOR2x1_ASAP7_75t_SL g986 ( .A(n_691), .B(n_539), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_791), .Y(n_987) );
INVxp33_ASAP7_75t_SL g988 ( .A(n_828), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_717), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_811), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_808), .B(n_16), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_719), .A2(n_539), .B1(n_566), .B2(n_553), .Y(n_992) );
INVxp67_ASAP7_75t_L g993 ( .A(n_785), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_809), .B(n_17), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_726), .A2(n_539), .B1(n_590), .B2(n_567), .C(n_580), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_689), .B(n_17), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_897), .B(n_689), .Y(n_997) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_878), .A2(n_739), .B1(n_732), .B2(n_742), .C(n_736), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_869), .A2(n_888), .B1(n_892), .B2(n_887), .C(n_952), .Y(n_999) );
BUFx6f_ASAP7_75t_L g1000 ( .A(n_936), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_859), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_869), .B(n_698), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_892), .A2(n_827), .B1(n_731), .B2(n_704), .C(n_698), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_958), .A2(n_781), .B1(n_695), .B2(n_799), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_937), .B(n_704), .Y(n_1005) );
OA21x2_ASAP7_75t_L g1006 ( .A1(n_834), .A2(n_567), .B(n_566), .Y(n_1006) );
BUFx2_ASAP7_75t_L g1007 ( .A(n_931), .Y(n_1007) );
AND2x4_ASAP7_75t_L g1008 ( .A(n_889), .B(n_691), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_929), .B(n_785), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_988), .A2(n_799), .B1(n_815), .B2(n_816), .Y(n_1010) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_897), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_975), .A2(n_815), .B1(n_731), .B2(n_768), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_871), .Y(n_1013) );
INVx8_ASAP7_75t_L g1014 ( .A(n_879), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_874), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_933), .B(n_823), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_848), .A2(n_762), .B1(n_765), .B2(n_728), .C(n_801), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_975), .A2(n_728), .B1(n_782), .B2(n_768), .Y(n_1018) );
OAI211xp5_ASAP7_75t_SL g1019 ( .A1(n_854), .A2(n_796), .B(n_801), .C(n_782), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_850), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_948), .B(n_796), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_979), .A2(n_831), .B1(n_778), .B2(n_716), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_972), .A2(n_932), .B1(n_955), .B2(n_976), .Y(n_1023) );
OAI21x1_ASAP7_75t_L g1024 ( .A1(n_843), .A2(n_818), .B(n_567), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_881), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_897), .A2(n_812), .B1(n_765), .B2(n_762), .Y(n_1026) );
OAI211xp5_ASAP7_75t_L g1027 ( .A1(n_848), .A2(n_818), .B(n_716), .C(n_725), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_948), .B(n_884), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_979), .A2(n_831), .B1(n_778), .B2(n_716), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_939), .A2(n_716), .B1(n_725), .B2(n_812), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_876), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_858), .B(n_19), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_939), .A2(n_778), .B1(n_725), .B2(n_758), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_877), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_886), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_854), .A2(n_725), .B1(n_758), .B2(n_737), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_879), .A2(n_895), .B1(n_979), .B2(n_860), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1038 ( .A1(n_879), .A2(n_724), .B1(n_747), .B2(n_744), .Y(n_1038) );
OR2x6_ASAP7_75t_L g1039 ( .A(n_853), .B(n_724), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_895), .A2(n_747), .B1(n_760), .B2(n_744), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_916), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_913), .B(n_737), .Y(n_1042) );
AOI21xp33_ASAP7_75t_L g1043 ( .A1(n_947), .A2(n_760), .B(n_747), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1044 ( .A(n_853), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_950), .A2(n_760), .B1(n_747), .B2(n_758), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1046 ( .A1(n_962), .A2(n_760), .B1(n_777), .B2(n_737), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_840), .A2(n_777), .B1(n_539), .B2(n_570), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_956), .A2(n_777), .B1(n_539), .B2(n_590), .C(n_566), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_922), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_924), .A2(n_570), .B1(n_590), .B2(n_580), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_913), .B(n_19), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_835), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_851), .B(n_21), .Y(n_1053) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_908), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_846), .A2(n_570), .B1(n_590), .B2(n_580), .Y(n_1055) );
AO21x2_ASAP7_75t_L g1056 ( .A1(n_961), .A2(n_570), .B(n_563), .Y(n_1056) );
OAI21xp33_ASAP7_75t_L g1057 ( .A1(n_875), .A2(n_575), .B(n_563), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_866), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_938), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_954), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1060) );
AOI222xp33_ASAP7_75t_L g1061 ( .A1(n_880), .A2(n_22), .B1(n_23), .B2(n_24), .C1(n_25), .C2(n_26), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1062 ( .A1(n_971), .A2(n_29), .B1(n_26), .B2(n_27), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_950), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_891), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_922), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_857), .Y(n_1066) );
AO31x2_ASAP7_75t_L g1067 ( .A1(n_961), .A2(n_33), .A3(n_30), .B(n_32), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_918), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g1069 ( .A(n_936), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_918), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_991), .A2(n_575), .B1(n_586), .B2(n_563), .Y(n_1071) );
NAND4xp25_ASAP7_75t_L g1072 ( .A(n_956), .B(n_35), .C(n_32), .D(n_33), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_971), .A2(n_38), .B1(n_36), .B2(n_37), .Y(n_1073) );
OAI211xp5_ASAP7_75t_SL g1074 ( .A1(n_912), .A2(n_41), .B(n_38), .C(n_40), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_902), .Y(n_1075) );
AOI222xp33_ASAP7_75t_L g1076 ( .A1(n_841), .A2(n_40), .B1(n_42), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_857), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_836), .B(n_42), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1079 ( .A1(n_970), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_985), .A2(n_592), .B1(n_586), .B2(n_575), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_963), .Y(n_1081) );
INVx3_ASAP7_75t_L g1082 ( .A(n_889), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_974), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_842), .B(n_861), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_959), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_993), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_987), .A2(n_592), .B1(n_586), .B2(n_49), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_875), .A2(n_592), .B1(n_48), .B2(n_49), .C(n_50), .Y(n_1088) );
NAND2xp33_ASAP7_75t_R g1089 ( .A(n_927), .B(n_47), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_909), .A2(n_592), .B1(n_48), .B2(n_50), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_864), .A2(n_592), .B1(n_51), .B2(n_52), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_868), .Y(n_1092) );
AOI22x1_ASAP7_75t_L g1093 ( .A1(n_980), .A2(n_592), .B1(n_51), .B2(n_52), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_865), .A2(n_592), .B1(n_53), .B2(n_54), .Y(n_1094) );
OAI221xp5_ASAP7_75t_L g1095 ( .A1(n_905), .A2(n_592), .B1(n_55), .B2(n_56), .C(n_57), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_960), .A2(n_47), .B1(n_56), .B2(n_58), .Y(n_1096) );
AOI222xp33_ASAP7_75t_L g1097 ( .A1(n_935), .A2(n_59), .B1(n_60), .B2(n_61), .C1(n_62), .C2(n_63), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_855), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_868), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_906), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_915), .B(n_63), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_926), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_907), .A2(n_64), .B1(n_65), .B2(n_67), .Y(n_1103) );
INVx4_ASAP7_75t_L g1104 ( .A(n_921), .Y(n_1104) );
OAI21xp5_ASAP7_75t_L g1105 ( .A1(n_905), .A2(n_581), .B(n_67), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_982), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_994), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_907), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_849), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_928), .A2(n_72), .B1(n_73), .B2(n_75), .C(n_77), .Y(n_1110) );
BUFx3_ASAP7_75t_L g1111 ( .A(n_915), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_906), .Y(n_1112) );
OAI221xp5_ASAP7_75t_SL g1113 ( .A1(n_920), .A2(n_73), .B1(n_78), .B2(n_80), .C(n_81), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_882), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_940), .A2(n_78), .B1(n_80), .B2(n_81), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_946), .B(n_82), .Y(n_1116) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_990), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_944), .A2(n_83), .B1(n_84), .B2(n_85), .C(n_86), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_966), .B(n_83), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_919), .A2(n_84), .B1(n_85), .B2(n_87), .Y(n_1120) );
OR2x6_ASAP7_75t_L g1121 ( .A(n_890), .B(n_88), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_849), .A2(n_88), .B1(n_90), .B2(n_91), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_993), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g1124 ( .A(n_936), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_896), .B(n_90), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_910), .A2(n_91), .B1(n_92), .B2(n_94), .Y(n_1126) );
OAI211xp5_ASAP7_75t_L g1127 ( .A1(n_953), .A2(n_581), .B(n_94), .C(n_97), .Y(n_1127) );
INVxp67_ASAP7_75t_L g1128 ( .A(n_957), .Y(n_1128) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_945), .A2(n_581), .B(n_130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_893), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_896), .A2(n_92), .B1(n_98), .B2(n_99), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_867), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_1132) );
OAI22x1_ASAP7_75t_L g1133 ( .A1(n_941), .A2(n_100), .B1(n_102), .B2(n_103), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_957), .A2(n_102), .B1(n_103), .B2(n_104), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_943), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_863), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_1136) );
AOI221x1_ASAP7_75t_SL g1137 ( .A1(n_919), .A2(n_105), .B1(n_107), .B2(n_108), .C(n_109), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_911), .A2(n_109), .B1(n_110), .B2(n_113), .Y(n_1138) );
NAND2x1p5_ASAP7_75t_L g1139 ( .A(n_890), .B(n_110), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_911), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_1140) );
NAND2xp5_ASAP7_75t_SL g1141 ( .A(n_870), .B(n_581), .Y(n_1141) );
AO22x1_ASAP7_75t_L g1142 ( .A1(n_894), .A2(n_114), .B1(n_115), .B2(n_117), .Y(n_1142) );
INVx4_ASAP7_75t_L g1143 ( .A(n_921), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_904), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1145 ( .A(n_923), .B(n_118), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1049), .B(n_941), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1147 ( .A1(n_999), .A2(n_930), .B1(n_920), .B2(n_844), .C(n_856), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1049), .B(n_873), .Y(n_1148) );
AOI222xp33_ASAP7_75t_L g1149 ( .A1(n_1037), .A2(n_900), .B1(n_883), .B2(n_965), .C1(n_862), .C2(n_856), .Y(n_1149) );
AOI33xp33_ASAP7_75t_L g1150 ( .A1(n_1023), .A2(n_862), .A3(n_863), .B1(n_872), .B2(n_969), .B3(n_844), .Y(n_1150) );
AOI221xp5_ASAP7_75t_L g1151 ( .A1(n_1062), .A2(n_984), .B1(n_872), .B2(n_967), .C(n_847), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1041), .Y(n_1152) );
OAI211xp5_ASAP7_75t_SL g1153 ( .A1(n_1076), .A2(n_968), .B(n_969), .C(n_978), .Y(n_1153) );
OA21x2_ASAP7_75t_L g1154 ( .A1(n_1024), .A2(n_977), .B(n_981), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_1014), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_1072), .A2(n_943), .B1(n_996), .B2(n_845), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_1086), .Y(n_1157) );
OA21x2_ASAP7_75t_L g1158 ( .A1(n_1071), .A2(n_977), .B(n_981), .Y(n_1158) );
AOI33xp33_ASAP7_75t_L g1159 ( .A1(n_1023), .A2(n_845), .A3(n_989), .B1(n_942), .B2(n_934), .B3(n_901), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_1137), .A2(n_885), .B1(n_992), .B2(n_995), .C(n_903), .Y(n_1160) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_1022), .A2(n_925), .B(n_917), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_1062), .A2(n_885), .B1(n_899), .B2(n_852), .C(n_917), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g1163 ( .A1(n_1073), .A2(n_852), .B1(n_838), .B2(n_983), .C(n_992), .Y(n_1163) );
INVxp67_ASAP7_75t_R g1164 ( .A(n_1133), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1014), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1066), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_1074), .A2(n_894), .B1(n_983), .B2(n_838), .Y(n_1167) );
OAI221xp5_ASAP7_75t_L g1168 ( .A1(n_1128), .A2(n_973), .B1(n_964), .B2(n_898), .C(n_914), .Y(n_1168) );
NAND4xp25_ASAP7_75t_L g1169 ( .A(n_1097), .B(n_119), .C(n_120), .D(n_121), .Y(n_1169) );
AOI211xp5_ASAP7_75t_L g1170 ( .A1(n_1073), .A2(n_973), .B(n_964), .C(n_914), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_1022), .Y(n_1171) );
OAI31xp33_ASAP7_75t_L g1172 ( .A1(n_1120), .A2(n_949), .A3(n_951), .B(n_894), .Y(n_1172) );
AND2x4_ASAP7_75t_SL g1173 ( .A(n_1121), .B(n_936), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_1121), .A2(n_949), .B1(n_894), .B2(n_839), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1032), .B(n_121), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_1120), .A2(n_1121), .B1(n_1075), .B2(n_1064), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1086), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1065), .B(n_122), .Y(n_1178) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1077), .Y(n_1179) );
OA21x2_ASAP7_75t_L g1180 ( .A1(n_1071), .A2(n_833), .B(n_837), .Y(n_1180) );
AND2x4_ASAP7_75t_L g1181 ( .A(n_1082), .B(n_986), .Y(n_1181) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_1014), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1013), .Y(n_1183) );
OAI33xp33_ASAP7_75t_L g1184 ( .A1(n_1102), .A2(n_123), .A3(n_833), .B1(n_837), .B2(n_894), .B3(n_134), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1065), .B(n_123), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1111), .B(n_833), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1015), .Y(n_1187) );
OAI31xp33_ASAP7_75t_L g1188 ( .A1(n_1102), .A2(n_833), .A3(n_839), .B(n_837), .Y(n_1188) );
OAI211xp5_ASAP7_75t_SL g1189 ( .A1(n_1107), .A2(n_837), .B(n_132), .C(n_133), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1025), .Y(n_1190) );
NAND4xp25_ASAP7_75t_L g1191 ( .A(n_1089), .B(n_1061), .C(n_1145), .D(n_1134), .Y(n_1191) );
OAI31xp33_ASAP7_75t_L g1192 ( .A1(n_1079), .A2(n_839), .A3(n_140), .B(n_142), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_1110), .A2(n_839), .B1(n_581), .B2(n_144), .Y(n_1193) );
AOI211xp5_ASAP7_75t_L g1194 ( .A1(n_1079), .A2(n_129), .B(n_143), .C(n_145), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1035), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1113), .A2(n_581), .B1(n_149), .B2(n_150), .C(n_151), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1020), .B(n_148), .Y(n_1197) );
AOI33xp33_ASAP7_75t_L g1198 ( .A1(n_1096), .A2(n_153), .A3(n_154), .B1(n_155), .B2(n_156), .B3(n_157), .Y(n_1198) );
OAI22xp33_ASAP7_75t_L g1199 ( .A1(n_1139), .A2(n_158), .B1(n_160), .B2(n_164), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1034), .B(n_167), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_1029), .A2(n_581), .B1(n_169), .B2(n_170), .Y(n_1201) );
OAI321xp33_ASAP7_75t_L g1202 ( .A1(n_1105), .A2(n_168), .A3(n_171), .B1(n_172), .B2(n_173), .C(n_174), .Y(n_1202) );
NOR3xp33_ASAP7_75t_L g1203 ( .A(n_1118), .B(n_175), .C(n_176), .Y(n_1203) );
OA21x2_ASAP7_75t_L g1204 ( .A1(n_1080), .A2(n_177), .B(n_178), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1101), .B(n_179), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1206 ( .A1(n_1139), .A2(n_180), .B1(n_184), .B2(n_185), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1028), .B(n_186), .Y(n_1207) );
OA21x2_ASAP7_75t_L g1208 ( .A1(n_1080), .A2(n_187), .B(n_188), .Y(n_1208) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_1117), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1011), .B(n_192), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g1211 ( .A1(n_1058), .A2(n_581), .B1(n_197), .B2(n_200), .C(n_208), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1095), .A2(n_581), .B1(n_209), .B2(n_210), .C(n_211), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1092), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1123), .B(n_196), .Y(n_1214) );
CKINVDCx20_ASAP7_75t_R g1215 ( .A(n_1001), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_1012), .A2(n_212), .B1(n_213), .B2(n_214), .C(n_215), .Y(n_1216) );
AOI22xp33_ASAP7_75t_SL g1217 ( .A1(n_1045), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_1051), .A2(n_220), .B1(n_221), .B2(n_222), .Y(n_1218) );
OAI221xp5_ASAP7_75t_L g1219 ( .A1(n_1012), .A2(n_223), .B1(n_224), .B2(n_228), .C(n_229), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1031), .Y(n_1220) );
AOI22xp33_ASAP7_75t_SL g1221 ( .A1(n_1093), .A2(n_1123), .B1(n_1135), .B2(n_1027), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1081), .B(n_230), .Y(n_1222) );
OAI31xp33_ASAP7_75t_L g1223 ( .A1(n_1029), .A2(n_233), .A3(n_234), .B(n_235), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g1224 ( .A1(n_1132), .A2(n_236), .B(n_241), .C(n_242), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_1126), .A2(n_243), .B1(n_244), .B2(n_249), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1054), .B(n_252), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1227 ( .A(n_1002), .B(n_253), .Y(n_1227) );
OAI221xp5_ASAP7_75t_SL g1228 ( .A1(n_1126), .A2(n_254), .B1(n_256), .B2(n_258), .C(n_259), .Y(n_1228) );
AOI33xp33_ASAP7_75t_L g1229 ( .A1(n_1096), .A2(n_268), .A3(n_272), .B1(n_274), .B2(n_275), .B3(n_277), .Y(n_1229) );
AOI21xp5_ASAP7_75t_L g1230 ( .A1(n_1057), .A2(n_278), .B(n_279), .Y(n_1230) );
AOI33xp33_ASAP7_75t_L g1231 ( .A1(n_1115), .A2(n_337), .A3(n_281), .B1(n_283), .B2(n_284), .B3(n_289), .Y(n_1231) );
OAI221xp5_ASAP7_75t_SL g1232 ( .A1(n_1115), .A2(n_280), .B1(n_291), .B2(n_292), .C(n_294), .Y(n_1232) );
OAI211xp5_ASAP7_75t_L g1233 ( .A1(n_1131), .A2(n_295), .B(n_296), .C(n_297), .Y(n_1233) );
NOR3xp33_ASAP7_75t_L g1234 ( .A(n_1125), .B(n_300), .C(n_302), .Y(n_1234) );
OAI31xp33_ASAP7_75t_L g1235 ( .A1(n_1019), .A2(n_304), .A3(n_305), .B(n_306), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_1109), .A2(n_308), .B1(n_314), .B2(n_316), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1000), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1007), .B(n_336), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1239 ( .A(n_1138), .B(n_319), .C(n_320), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1000), .Y(n_1240) );
OAI211xp5_ASAP7_75t_SL g1241 ( .A1(n_1085), .A2(n_326), .B(n_329), .C(n_330), .Y(n_1241) );
NOR2x1_ASAP7_75t_L g1242 ( .A(n_1104), .B(n_332), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1052), .B(n_333), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1083), .Y(n_1244) );
INVx1_ASAP7_75t_SL g1245 ( .A(n_1044), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1030), .A2(n_335), .B1(n_1033), .B2(n_1018), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1104), .B(n_1143), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_997), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1099), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1018), .A2(n_1090), .B1(n_1036), .B2(n_1010), .Y(n_1250) );
INVx5_ASAP7_75t_L g1251 ( .A(n_1039), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1090), .A2(n_1010), .B1(n_1063), .B2(n_1070), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_1068), .A2(n_1026), .B1(n_1094), .B2(n_1108), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1130), .B(n_1106), .Y(n_1254) );
OAI211xp5_ASAP7_75t_SL g1255 ( .A1(n_1140), .A2(n_1144), .B(n_1119), .C(n_1116), .Y(n_1255) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_1103), .A2(n_1108), .B1(n_1094), .B2(n_1003), .C(n_1127), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1114), .B(n_1143), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1103), .B(n_1112), .Y(n_1258) );
NAND4xp25_ASAP7_75t_L g1259 ( .A(n_1053), .B(n_1078), .C(n_1091), .D(n_1004), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_1088), .A2(n_1087), .B1(n_998), .B2(n_1004), .C(n_1098), .Y(n_1260) );
AOI21xp5_ASAP7_75t_L g1261 ( .A1(n_1038), .A2(n_1040), .B(n_1129), .Y(n_1261) );
AOI221xp5_ASAP7_75t_L g1262 ( .A1(n_1169), .A2(n_1122), .B1(n_1136), .B2(n_1142), .C(n_1084), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1186), .B(n_1100), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1166), .B(n_1067), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1183), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1157), .B(n_1177), .Y(n_1266) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1181), .B(n_1067), .Y(n_1267) );
OAI22xp33_ASAP7_75t_L g1268 ( .A1(n_1191), .A2(n_1046), .B1(n_1017), .B2(n_1082), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1187), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1254), .Y(n_1270) );
NAND4xp25_ASAP7_75t_L g1271 ( .A(n_1176), .B(n_1087), .C(n_1055), .D(n_1060), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1179), .B(n_1067), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1152), .B(n_1067), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1190), .B(n_1009), .Y(n_1274) );
INVx3_ASAP7_75t_L g1275 ( .A(n_1173), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1213), .B(n_1056), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1176), .A2(n_1149), .B1(n_1156), .B2(n_1172), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1195), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1249), .B(n_1056), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1180), .Y(n_1280) );
NAND3xp33_ASAP7_75t_L g1281 ( .A(n_1221), .B(n_1047), .C(n_1043), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_1156), .A2(n_1042), .B1(n_1021), .B2(n_1141), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_1259), .A2(n_1039), .B1(n_1048), .B2(n_1038), .Y(n_1283) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_1171), .A2(n_1008), .B1(n_1006), .B2(n_1039), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1244), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1157), .B(n_1006), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1287 ( .A(n_1165), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1220), .B(n_1005), .Y(n_1288) );
AND2x4_ASAP7_75t_L g1289 ( .A(n_1181), .B(n_1000), .Y(n_1289) );
OAI22xp33_ASAP7_75t_L g1290 ( .A1(n_1164), .A2(n_1016), .B1(n_1006), .B2(n_1008), .Y(n_1290) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1180), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1177), .B(n_1000), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1178), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1180), .B(n_1069), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1185), .Y(n_1295) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_1167), .A2(n_1050), .B1(n_1059), .B2(n_1069), .C(n_1124), .Y(n_1296) );
OAI221xp5_ASAP7_75t_L g1297 ( .A1(n_1167), .A2(n_1069), .B1(n_1124), .B2(n_1260), .C(n_1209), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1257), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1146), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1300 ( .A(n_1247), .Y(n_1300) );
OR2x6_ASAP7_75t_L g1301 ( .A(n_1174), .B(n_1069), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1148), .B(n_1124), .Y(n_1302) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1237), .Y(n_1303) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1237), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1258), .B(n_1124), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1240), .B(n_1159), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1247), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1226), .Y(n_1308) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1240), .Y(n_1309) );
OAI33xp33_ASAP7_75t_L g1310 ( .A1(n_1238), .A2(n_1199), .A3(n_1206), .B1(n_1250), .B2(n_1255), .B3(n_1248), .Y(n_1310) );
NOR3xp33_ASAP7_75t_SL g1311 ( .A(n_1210), .B(n_1206), .C(n_1199), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_1147), .A2(n_1153), .B1(n_1256), .B2(n_1253), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_1252), .A2(n_1203), .B1(n_1151), .B2(n_1175), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1314 ( .A1(n_1170), .A2(n_1193), .B1(n_1194), .B2(n_1225), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1159), .B(n_1188), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1173), .B(n_1214), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_1193), .A2(n_1225), .B1(n_1228), .B2(n_1232), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1242), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1150), .B(n_1155), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1204), .Y(n_1320) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1154), .Y(n_1321) );
BUFx2_ASAP7_75t_L g1322 ( .A(n_1251), .Y(n_1322) );
OAI31xp33_ASAP7_75t_L g1323 ( .A1(n_1210), .A2(n_1192), .A3(n_1182), .B(n_1224), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1150), .B(n_1165), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_1236), .A2(n_1196), .B1(n_1160), .B2(n_1163), .Y(n_1325) );
INVx4_ASAP7_75t_L g1326 ( .A(n_1251), .Y(n_1326) );
INVx1_ASAP7_75t_SL g1327 ( .A(n_1245), .Y(n_1327) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1154), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_1184), .A2(n_1227), .B1(n_1212), .B2(n_1246), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1207), .B(n_1205), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1243), .B(n_1227), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1162), .B(n_1251), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1333 ( .A1(n_1236), .A2(n_1251), .B1(n_1218), .B2(n_1216), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1158), .B(n_1200), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_1189), .A2(n_1222), .B1(n_1161), .B2(n_1211), .C(n_1202), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1197), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1231), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1231), .B(n_1198), .Y(n_1338) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_1234), .A2(n_1201), .B1(n_1215), .B2(n_1239), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1340 ( .A(n_1204), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1158), .B(n_1204), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1208), .Y(n_1342) );
OAI33xp33_ASAP7_75t_L g1343 ( .A1(n_1241), .A2(n_1229), .A3(n_1198), .B1(n_1223), .B2(n_1235), .B3(n_1233), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1344 ( .A1(n_1261), .A2(n_1208), .B(n_1230), .Y(n_1344) );
AOI33xp33_ASAP7_75t_L g1345 ( .A1(n_1218), .A2(n_1217), .A3(n_1229), .B1(n_1219), .B2(n_1208), .B3(n_1158), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1154), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1168), .Y(n_1347) );
NAND2x1p5_ASAP7_75t_L g1348 ( .A(n_1181), .B(n_1251), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1186), .Y(n_1349) );
NOR4xp25_ASAP7_75t_L g1350 ( .A(n_1327), .B(n_1277), .C(n_1312), .D(n_1278), .Y(n_1350) );
INVxp67_ASAP7_75t_L g1351 ( .A(n_1300), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1265), .Y(n_1352) );
INVxp67_ASAP7_75t_L g1353 ( .A(n_1287), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1265), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1269), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1349), .B(n_1305), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1269), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1310), .A2(n_1313), .B1(n_1325), .B2(n_1262), .Y(n_1358) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_1267), .B(n_1305), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1280), .Y(n_1360) );
INVx2_ASAP7_75t_SL g1361 ( .A(n_1322), .Y(n_1361) );
OAI332xp33_ASAP7_75t_L g1362 ( .A1(n_1270), .A2(n_1268), .A3(n_1319), .B1(n_1293), .B2(n_1295), .B3(n_1274), .C1(n_1299), .C2(n_1324), .Y(n_1362) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_1266), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1349), .B(n_1266), .Y(n_1364) );
NOR3xp33_ASAP7_75t_SL g1365 ( .A(n_1323), .B(n_1343), .C(n_1314), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1298), .B(n_1285), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1285), .B(n_1307), .Y(n_1367) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_1318), .B(n_1281), .C(n_1297), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1263), .B(n_1302), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1263), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1273), .B(n_1309), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1288), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1308), .B(n_1336), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1287), .B(n_1315), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1315), .B(n_1292), .Y(n_1375) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1303), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1334), .B(n_1264), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1334), .B(n_1264), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1303), .Y(n_1379) );
NOR3xp33_ASAP7_75t_L g1380 ( .A(n_1318), .B(n_1271), .C(n_1339), .Y(n_1380) );
INVxp67_ASAP7_75t_L g1381 ( .A(n_1292), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1272), .B(n_1276), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1383 ( .A(n_1267), .B(n_1294), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1384 ( .A1(n_1337), .A2(n_1306), .B1(n_1338), .B2(n_1290), .C(n_1317), .Y(n_1384) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_1330), .B(n_1331), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1304), .B(n_1309), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1304), .B(n_1272), .Y(n_1387) );
O2A1O1Ixp33_ASAP7_75t_L g1388 ( .A1(n_1330), .A2(n_1311), .B(n_1347), .C(n_1333), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1286), .Y(n_1389) );
OAI21xp5_ASAP7_75t_SL g1390 ( .A1(n_1348), .A2(n_1283), .B(n_1322), .Y(n_1390) );
INVx2_ASAP7_75t_SL g1391 ( .A(n_1348), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1276), .B(n_1279), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1286), .B(n_1346), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1316), .B(n_1348), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1306), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1279), .B(n_1267), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1282), .B(n_1347), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1316), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1291), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1275), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1275), .Y(n_1401) );
AND2x4_ASAP7_75t_L g1402 ( .A(n_1294), .B(n_1332), .Y(n_1402) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1321), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1275), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1341), .B(n_1346), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1296), .B(n_1332), .Y(n_1406) );
NOR3xp33_ASAP7_75t_SL g1407 ( .A(n_1335), .B(n_1344), .C(n_1342), .Y(n_1407) );
INVx2_ASAP7_75t_L g1408 ( .A(n_1321), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1341), .B(n_1328), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1326), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1328), .B(n_1320), .Y(n_1411) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1342), .Y(n_1412) );
NOR3xp33_ASAP7_75t_L g1413 ( .A(n_1345), .B(n_1326), .C(n_1284), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1326), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1367), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1363), .B(n_1289), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1352), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1372), .B(n_1289), .Y(n_1418) );
O2A1O1Ixp33_ASAP7_75t_L g1419 ( .A1(n_1365), .A2(n_1329), .B(n_1340), .C(n_1301), .Y(n_1419) );
AOI33xp33_ASAP7_75t_L g1420 ( .A1(n_1358), .A2(n_1289), .A3(n_1301), .B1(n_1340), .B2(n_1345), .B3(n_1350), .Y(n_1420) );
NAND2x1_ASAP7_75t_L g1421 ( .A(n_1391), .B(n_1301), .Y(n_1421) );
OR2x2_ASAP7_75t_L g1422 ( .A(n_1395), .B(n_1301), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_1374), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1366), .Y(n_1424) );
INVxp67_ASAP7_75t_L g1425 ( .A(n_1375), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1354), .Y(n_1426) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_1385), .B(n_1351), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1355), .Y(n_1428) );
INVxp67_ASAP7_75t_SL g1429 ( .A(n_1361), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1357), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1370), .B(n_1385), .Y(n_1431) );
NOR2xp33_ASAP7_75t_L g1432 ( .A(n_1362), .B(n_1373), .Y(n_1432) );
OR2x6_ASAP7_75t_L g1433 ( .A(n_1390), .B(n_1391), .Y(n_1433) );
AOI21xp5_ASAP7_75t_L g1434 ( .A1(n_1388), .A2(n_1413), .B(n_1361), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1377), .B(n_1378), .Y(n_1435) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_1383), .B(n_1359), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1364), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1412), .Y(n_1438) );
NOR3xp33_ASAP7_75t_SL g1439 ( .A(n_1384), .B(n_1397), .C(n_1406), .Y(n_1439) );
BUFx3_ASAP7_75t_L g1440 ( .A(n_1410), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1364), .B(n_1393), .Y(n_1441) );
AOI321xp33_ASAP7_75t_L g1442 ( .A1(n_1358), .A2(n_1380), .A3(n_1406), .B1(n_1368), .B2(n_1398), .C(n_1356), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1356), .Y(n_1443) );
OA211x2_ASAP7_75t_L g1444 ( .A1(n_1353), .A2(n_1381), .B(n_1407), .C(n_1394), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1382), .B(n_1392), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1393), .B(n_1389), .Y(n_1446) );
INVx2_ASAP7_75t_L g1447 ( .A(n_1412), .Y(n_1447) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1360), .Y(n_1448) );
BUFx2_ASAP7_75t_L g1449 ( .A(n_1383), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1382), .B(n_1392), .Y(n_1450) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1360), .Y(n_1451) );
NAND2x1p5_ASAP7_75t_L g1452 ( .A(n_1414), .B(n_1404), .Y(n_1452) );
NOR2x1_ASAP7_75t_L g1453 ( .A(n_1400), .B(n_1401), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1371), .B(n_1369), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1371), .Y(n_1455) );
HB1xp67_ASAP7_75t_L g1456 ( .A(n_1386), .Y(n_1456) );
INVxp67_ASAP7_75t_L g1457 ( .A(n_1386), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1396), .B(n_1405), .Y(n_1458) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_1432), .A2(n_1402), .B1(n_1359), .B2(n_1396), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_1433), .A2(n_1383), .B1(n_1402), .B2(n_1359), .Y(n_1460) );
INVxp67_ASAP7_75t_SL g1461 ( .A(n_1456), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1438), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1438), .Y(n_1463) );
XNOR2xp5_ASAP7_75t_L g1464 ( .A(n_1439), .B(n_1402), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1417), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1466 ( .A(n_1457), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1435), .B(n_1409), .Y(n_1467) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1417), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1435), .B(n_1409), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1455), .B(n_1411), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1455), .B(n_1411), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1415), .B(n_1376), .Y(n_1472) );
OAI21xp33_ASAP7_75t_SL g1473 ( .A1(n_1433), .A2(n_1379), .B(n_1387), .Y(n_1473) );
A2O1A1Ixp33_ASAP7_75t_SL g1474 ( .A1(n_1419), .A2(n_1399), .B(n_1403), .C(n_1408), .Y(n_1474) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_1433), .A2(n_1387), .B1(n_1403), .B2(n_1408), .Y(n_1475) );
AND3x2_ASAP7_75t_L g1476 ( .A(n_1429), .B(n_1449), .C(n_1420), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1424), .B(n_1437), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1426), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1426), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1458), .B(n_1450), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1458), .B(n_1450), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1445), .B(n_1443), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1445), .B(n_1449), .Y(n_1483) );
XNOR2x2_ASAP7_75t_L g1484 ( .A(n_1434), .B(n_1453), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1428), .Y(n_1485) );
A2O1A1Ixp33_ASAP7_75t_SL g1486 ( .A1(n_1423), .A2(n_1425), .B(n_1427), .C(n_1416), .Y(n_1486) );
XNOR2x1_ASAP7_75t_L g1487 ( .A(n_1431), .B(n_1444), .Y(n_1487) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1428), .Y(n_1488) );
AND2x4_ASAP7_75t_SL g1489 ( .A(n_1436), .B(n_1433), .Y(n_1489) );
AOI211xp5_ASAP7_75t_L g1490 ( .A1(n_1436), .A2(n_1422), .B(n_1441), .C(n_1418), .Y(n_1490) );
INVxp67_ASAP7_75t_L g1491 ( .A(n_1440), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1454), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1454), .Y(n_1493) );
HB1xp67_ASAP7_75t_L g1494 ( .A(n_1446), .Y(n_1494) );
NOR2xp33_ASAP7_75t_L g1495 ( .A(n_1446), .B(n_1436), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1447), .B(n_1422), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1430), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1447), .B(n_1448), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1430), .Y(n_1499) );
AOI21xp5_ASAP7_75t_L g1500 ( .A1(n_1421), .A2(n_1452), .B(n_1440), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1448), .B(n_1451), .Y(n_1501) );
INVx1_ASAP7_75t_SL g1502 ( .A(n_1421), .Y(n_1502) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_1442), .A2(n_1380), .B1(n_1365), .B2(n_1432), .Y(n_1503) );
NAND2xp33_ASAP7_75t_SL g1504 ( .A(n_1451), .B(n_1452), .Y(n_1504) );
INVxp67_ASAP7_75t_SL g1505 ( .A(n_1452), .Y(n_1505) );
AOI22xp5_ASAP7_75t_L g1506 ( .A1(n_1432), .A2(n_1380), .B1(n_1365), .B2(n_1358), .Y(n_1506) );
INVx2_ASAP7_75t_L g1507 ( .A(n_1483), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_1464), .A2(n_1489), .B1(n_1487), .B2(n_1490), .Y(n_1508) );
AOI221xp5_ASAP7_75t_L g1509 ( .A1(n_1503), .A2(n_1506), .B1(n_1486), .B2(n_1464), .C(n_1466), .Y(n_1509) );
AOI321xp33_ASAP7_75t_L g1510 ( .A1(n_1460), .A2(n_1475), .A3(n_1459), .B1(n_1461), .B2(n_1483), .C(n_1495), .Y(n_1510) );
AOI21xp33_ASAP7_75t_SL g1511 ( .A1(n_1487), .A2(n_1473), .B(n_1460), .Y(n_1511) );
NAND2xp5_ASAP7_75t_SL g1512 ( .A(n_1473), .B(n_1489), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1466), .Y(n_1513) );
XNOR2xp5_ASAP7_75t_L g1514 ( .A(n_1459), .B(n_1476), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1480), .B(n_1481), .Y(n_1515) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_1476), .A2(n_1475), .B1(n_1492), .B2(n_1493), .Y(n_1516) );
NAND2x1_ASAP7_75t_SL g1517 ( .A(n_1494), .B(n_1484), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1480), .B(n_1481), .Y(n_1518) );
AOI21xp33_ASAP7_75t_SL g1519 ( .A1(n_1491), .A2(n_1484), .B(n_1486), .Y(n_1519) );
O2A1O1Ixp33_ASAP7_75t_L g1520 ( .A1(n_1474), .A2(n_1461), .B(n_1500), .C(n_1505), .Y(n_1520) );
NAND2xp33_ASAP7_75t_SL g1521 ( .A(n_1469), .B(n_1467), .Y(n_1521) );
AOI21xp5_ASAP7_75t_L g1522 ( .A1(n_1512), .A2(n_1504), .B(n_1502), .Y(n_1522) );
A2O1A1Ixp33_ASAP7_75t_SL g1523 ( .A1(n_1520), .A2(n_1478), .B(n_1488), .C(n_1468), .Y(n_1523) );
AOI221xp5_ASAP7_75t_L g1524 ( .A1(n_1509), .A2(n_1511), .B1(n_1508), .B2(n_1519), .C(n_1514), .Y(n_1524) );
XNOR2x1_ASAP7_75t_L g1525 ( .A(n_1516), .B(n_1482), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1526 ( .A(n_1513), .B(n_1482), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_1521), .A2(n_1477), .B1(n_1504), .B2(n_1472), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1518), .Y(n_1528) );
AOI211xp5_ASAP7_75t_SL g1529 ( .A1(n_1517), .A2(n_1470), .B(n_1471), .C(n_1469), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1507), .Y(n_1530) );
AOI21xp5_ASAP7_75t_L g1531 ( .A1(n_1520), .A2(n_1471), .B(n_1470), .Y(n_1531) );
NOR4xp25_ASAP7_75t_L g1532 ( .A(n_1524), .B(n_1510), .C(n_1515), .D(n_1467), .Y(n_1532) );
NOR3xp33_ASAP7_75t_SL g1533 ( .A(n_1522), .B(n_1501), .C(n_1478), .Y(n_1533) );
OAI211xp5_ASAP7_75t_SL g1534 ( .A1(n_1529), .A2(n_1499), .B(n_1497), .C(n_1465), .Y(n_1534) );
OAI22xp5_ASAP7_75t_SL g1535 ( .A1(n_1527), .A2(n_1468), .B1(n_1479), .B2(n_1465), .Y(n_1535) );
AOI22xp5_ASAP7_75t_L g1536 ( .A1(n_1525), .A2(n_1496), .B1(n_1479), .B2(n_1488), .Y(n_1536) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1528), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1537), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_1536), .A2(n_1527), .B1(n_1531), .B2(n_1526), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1535), .Y(n_1540) );
NOR2xp33_ASAP7_75t_L g1541 ( .A(n_1534), .B(n_1530), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1538), .Y(n_1542) );
OAI221xp5_ASAP7_75t_L g1543 ( .A1(n_1540), .A2(n_1532), .B1(n_1523), .B2(n_1533), .C(n_1485), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1541), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1542), .Y(n_1545) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1542), .Y(n_1546) );
INVxp67_ASAP7_75t_SL g1547 ( .A(n_1546), .Y(n_1547) );
AO21x1_ASAP7_75t_L g1548 ( .A1(n_1545), .A2(n_1544), .B(n_1539), .Y(n_1548) );
OAI21x1_ASAP7_75t_SL g1549 ( .A1(n_1548), .A2(n_1543), .B(n_1485), .Y(n_1549) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_1549), .A2(n_1547), .B1(n_1462), .B2(n_1463), .C(n_1498), .Y(n_1550) );
endmodule