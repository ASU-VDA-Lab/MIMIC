module fake_jpeg_9314_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVxp67_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_19),
.Y(n_23)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_18)
);

A2O1A1O1Ixp25_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_8),
.B(n_5),
.C(n_6),
.D(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_3),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_12),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_17),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_7),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_4),
.C(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_37),
.B(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_38),
.C(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_41),
.A3(n_46),
.B1(n_45),
.B2(n_31),
.C1(n_39),
.C2(n_22),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.C(n_48),
.Y(n_50)
);


endmodule