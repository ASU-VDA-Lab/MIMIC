module fake_netlist_6_4268_n_31 (n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_31);

input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_31;

wire n_16;
wire n_9;
wire n_8;
wire n_18;
wire n_21;
wire n_10;
wire n_24;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_7;
wire n_30;
wire n_19;
wire n_29;
wire n_25;

INVx2_ASAP7_75t_SL g7 ( 
.A(n_3),
.Y(n_7)
);

AND2x4_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_4),
.Y(n_8)
);

OAI21x1_ASAP7_75t_L g9 ( 
.A1(n_4),
.A2(n_5),
.B(n_3),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_8),
.B(n_7),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_15),
.Y(n_17)
);

OA21x2_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_9),
.B(n_12),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_8),
.A3(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR3xp33_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_25),
.C(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_11),
.B1(n_8),
.B2(n_18),
.Y(n_29)
);

AO21x2_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_23),
.B(n_18),
.Y(n_30)
);

AO221x2_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_2),
.B1(n_10),
.B2(n_23),
.C(n_28),
.Y(n_31)
);


endmodule