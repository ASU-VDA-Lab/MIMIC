module fake_netlist_1_1124_n_994 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_994);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_994;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_627;
wire n_532;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_158), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_138), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_100), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_12), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_72), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_78), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_133), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_71), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_123), .Y(n_252) );
INVxp33_ASAP7_75t_SL g253 ( .A(n_120), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_225), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_99), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_184), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_10), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_2), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_70), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_31), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_48), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_238), .Y(n_262) );
CKINVDCx14_ASAP7_75t_R g263 ( .A(n_194), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_193), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_171), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_156), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_17), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_73), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_231), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_68), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_19), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_163), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_39), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_46), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_85), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
BUFx5_ASAP7_75t_L g277 ( .A(n_203), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_112), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_154), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_137), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_79), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_223), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_16), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_83), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_61), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_200), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_131), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_86), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_52), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_98), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_81), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_179), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_48), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_20), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_125), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_149), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_66), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_59), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_1), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_30), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_132), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_197), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_130), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_172), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_28), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_232), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_229), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_122), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_114), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_185), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_49), .Y(n_313) );
INVxp33_ASAP7_75t_L g314 ( .A(n_118), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_19), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_169), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_103), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_23), .Y(n_318) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_212), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_214), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_190), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_215), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_95), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_25), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_90), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_146), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_167), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_17), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_195), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_29), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_205), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_128), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_111), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_208), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_126), .Y(n_335) );
CKINVDCx16_ASAP7_75t_R g336 ( .A(n_39), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_75), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_102), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_27), .B(n_202), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_84), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_54), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_110), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_209), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_143), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_136), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_192), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_25), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_217), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_80), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_162), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_177), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_213), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_54), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_104), .Y(n_354) );
INVxp33_ASAP7_75t_SL g355 ( .A(n_106), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_181), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_175), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_189), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_121), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_60), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_166), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_115), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_124), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_52), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_91), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_77), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_92), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_8), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_107), .Y(n_369) );
XNOR2xp5_ASAP7_75t_L g370 ( .A(n_16), .B(n_127), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_165), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_174), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_237), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_40), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_152), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_36), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_5), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_277), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_257), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_314), .B(n_0), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_257), .B(n_0), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_336), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_274), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_314), .B(n_1), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_248), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_277), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_251), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_315), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_277), .Y(n_389) );
NOR2xp33_ASAP7_75t_R g390 ( .A(n_263), .B(n_63), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_246), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_258), .B(n_2), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_315), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_277), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_274), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_262), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_244), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_277), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_293), .B(n_3), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_247), .B(n_3), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_245), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_263), .B(n_4), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_261), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_277), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_249), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_262), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_250), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_277), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_399), .B(n_270), .Y(n_409) );
OR2x6_ASAP7_75t_L g410 ( .A(n_403), .B(n_319), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_403), .B(n_356), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_397), .B(n_292), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_397), .B(n_308), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_406), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_382), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_401), .B(n_337), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_381), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_401), .B(n_254), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_405), .B(n_254), .Y(n_422) );
AND2x6_ASAP7_75t_L g423 ( .A(n_399), .B(n_375), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_380), .B(n_261), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_402), .B(n_243), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_392), .B(n_285), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
BUFx8_ASAP7_75t_SL g430 ( .A(n_383), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_405), .B(n_287), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g433 ( .A(n_402), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_407), .B(n_287), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_388), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_399), .B(n_260), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_392), .B(n_267), .Y(n_444) );
INVx6_ASAP7_75t_L g445 ( .A(n_396), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_407), .B(n_299), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_392), .B(n_271), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_393), .B(n_299), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_448), .B(n_385), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_448), .B(n_387), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_427), .A2(n_269), .B1(n_331), .B2(n_272), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_451), .A2(n_272), .B1(n_331), .B2(n_269), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_427), .B(n_243), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_411), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_441), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_424), .B(n_378), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_429), .A2(n_386), .B1(n_389), .B2(n_378), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_442), .Y(n_463) );
AOI21x1_ASAP7_75t_L g464 ( .A1(n_421), .A2(n_386), .B(n_378), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_416), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_413), .A2(n_408), .B(n_389), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_433), .B(n_353), .C(n_290), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_432), .B(n_253), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_409), .B(n_266), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_435), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_450), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_410), .B(n_273), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_409), .B(n_266), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_439), .B(n_386), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_439), .B(n_389), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_412), .B(n_285), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
OAI21xp33_ASAP7_75t_SL g481 ( .A1(n_420), .A2(n_398), .B(n_394), .Y(n_481) );
AND2x6_ASAP7_75t_SL g482 ( .A(n_430), .B(n_395), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_425), .A2(n_346), .B1(n_324), .B2(n_328), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_414), .B(n_275), .Y(n_484) );
BUFx4f_ASAP7_75t_L g485 ( .A(n_410), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_414), .B(n_275), .Y(n_486) );
NAND2x2_ASAP7_75t_L g487 ( .A(n_418), .B(n_375), .Y(n_487) );
INVx5_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_415), .B(n_286), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_436), .A2(n_398), .B1(n_404), .B2(n_394), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_426), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_444), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_443), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_444), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_419), .B(n_322), .Y(n_497) );
NAND2xp33_ASAP7_75t_L g498 ( .A(n_423), .B(n_390), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_447), .A2(n_346), .B1(n_324), .B2(n_328), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_416), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_419), .B(n_322), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_447), .B(n_394), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_438), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_449), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_421), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_434), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_446), .B(n_345), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_434), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_434), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_422), .B(n_398), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_422), .B(n_253), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_431), .B(n_345), .Y(n_512) );
INVx5_ASAP7_75t_L g513 ( .A(n_434), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_431), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_440), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_440), .B(n_355), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_440), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_440), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_451), .B(n_404), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_448), .B(n_355), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_427), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_424), .A2(n_408), .B1(n_404), .B2(n_296), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_418), .A2(n_360), .B1(n_370), .B2(n_341), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_416), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_451), .B(n_408), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_451), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_435), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_528), .A2(n_360), .B1(n_368), .B2(n_313), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_477), .B(n_350), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_458), .A2(n_295), .B1(n_301), .B2(n_300), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_492), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_454), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_480), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_521), .A2(n_264), .B1(n_318), .B2(n_307), .Y(n_537) );
OR2x6_ASAP7_75t_SL g538 ( .A(n_499), .B(n_350), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_471), .B(n_302), .Y(n_539) );
OR2x6_ASAP7_75t_L g540 ( .A(n_474), .B(n_496), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_521), .B(n_366), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_453), .B(n_339), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_476), .A2(n_362), .B(n_338), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_488), .B(n_366), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_480), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_492), .A2(n_330), .B(n_364), .C(n_347), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_458), .A2(n_374), .B1(n_377), .B2(n_376), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_485), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_493), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_476), .A2(n_255), .B(n_252), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_452), .B(n_298), .Y(n_552) );
INVx4_ASAP7_75t_SL g553 ( .A(n_524), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_520), .B(n_309), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_455), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_494), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_522), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_SL g558 ( .A1(n_468), .A2(n_391), .B(n_317), .C(n_343), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_479), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_468), .A2(n_283), .B1(n_246), .B2(n_396), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_478), .A2(n_259), .B(n_256), .Y(n_562) );
OR2x6_ASAP7_75t_L g563 ( .A(n_495), .B(n_246), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_483), .B(n_4), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_478), .A2(n_268), .B(n_265), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_504), .A2(n_523), .B1(n_473), .B2(n_459), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_491), .Y(n_567) );
NOR2xp67_ASAP7_75t_SL g568 ( .A(n_488), .B(n_371), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_519), .A2(n_278), .B(n_276), .Y(n_570) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_467), .B(n_246), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_503), .B(n_333), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g573 ( .A1(n_467), .A2(n_280), .B(n_281), .C(n_279), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_469), .A2(n_283), .B1(n_284), .B2(n_282), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_519), .A2(n_289), .B(n_288), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_452), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_475), .B(n_291), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_456), .B(n_294), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_457), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_488), .B(n_283), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_488), .Y(n_582) );
INVx4_ASAP7_75t_L g583 ( .A(n_513), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_507), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_527), .A2(n_297), .B1(n_304), .B2(n_303), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_481), .A2(n_310), .B(n_306), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_484), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_502), .B(n_311), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_502), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_527), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_472), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_511), .A2(n_283), .B1(n_396), .B2(n_406), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_486), .B(n_5), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_489), .A2(n_344), .B1(n_312), .B2(n_373), .C1(n_372), .C2(n_316), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_463), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_497), .B(n_320), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_517), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_513), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_464), .Y(n_600) );
O2A1O1Ixp5_ASAP7_75t_L g601 ( .A1(n_516), .A2(n_317), .B(n_343), .C(n_305), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_513), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_460), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_462), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_511), .A2(n_406), .B1(n_321), .B2(n_325), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_466), .A2(n_351), .B(n_323), .C(n_326), .Y(n_606) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_498), .B(n_327), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_501), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_514), .A2(n_406), .B1(n_354), .B2(n_352), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_460), .A2(n_510), .B(n_505), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_523), .B(n_329), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_510), .A2(n_334), .B(n_332), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g613 ( .A1(n_461), .A2(n_358), .B(n_335), .C(n_340), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_512), .B(n_6), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_461), .B(n_342), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_490), .B(n_6), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_490), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_513), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_525), .B(n_515), .Y(n_619) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_487), .B(n_348), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_487), .A2(n_406), .B1(n_363), .B2(n_361), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_470), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_462), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_462), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_470), .A2(n_365), .B1(n_367), .B2(n_357), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_518), .A2(n_359), .B(n_349), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_529), .B(n_7), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_529), .A2(n_369), .B1(n_349), .B2(n_305), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_508), .B(n_7), .Y(n_629) );
NOR2xp33_ASAP7_75t_SL g630 ( .A(n_465), .B(n_509), .Y(n_630) );
OR2x6_ASAP7_75t_L g631 ( .A(n_465), .B(n_391), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_509), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_509), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_SL g634 ( .A1(n_500), .A2(n_391), .B(n_117), .C(n_119), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_506), .B(n_8), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_509), .Y(n_636) );
INVx4_ASAP7_75t_L g637 ( .A(n_526), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_526), .B(n_9), .Y(n_638) );
CKINVDCx16_ASAP7_75t_R g639 ( .A(n_526), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_528), .B(n_391), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_528), .B(n_9), .Y(n_641) );
AO21x2_ASAP7_75t_L g642 ( .A1(n_600), .A2(n_65), .B(n_64), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_533), .B(n_11), .Y(n_643) );
AO31x2_ASAP7_75t_L g644 ( .A1(n_566), .A2(n_11), .A3(n_12), .B(n_13), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_617), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_604), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_616), .A2(n_14), .B1(n_15), .B2(n_18), .Y(n_647) );
AO21x2_ASAP7_75t_L g648 ( .A1(n_558), .A2(n_69), .B(n_67), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_639), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_540), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_579), .Y(n_651) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_566), .A2(n_606), .A3(n_613), .B(n_625), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_546), .A2(n_18), .B1(n_20), .B2(n_21), .C(n_22), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_559), .B(n_21), .Y(n_654) );
O2A1O1Ixp5_ASAP7_75t_L g655 ( .A1(n_601), .A2(n_140), .B(n_241), .C(n_240), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_576), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_656) );
OAI21x1_ASAP7_75t_L g657 ( .A1(n_636), .A2(n_76), .B(n_74), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_610), .A2(n_87), .B(n_82), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_530), .B(n_24), .Y(n_659) );
OAI21x1_ASAP7_75t_L g660 ( .A1(n_581), .A2(n_89), .B(n_88), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_592), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_550), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_581), .A2(n_94), .B(n_93), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_586), .A2(n_147), .B(n_239), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_596), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_596), .B(n_29), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_538), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_567), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_530), .B(n_32), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_534), .B(n_33), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_604), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_556), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_604), .Y(n_674) );
OA21x2_ASAP7_75t_L g675 ( .A1(n_586), .A2(n_153), .B(n_236), .Y(n_675) );
OR2x6_ASAP7_75t_L g676 ( .A(n_540), .B(n_34), .Y(n_676) );
AO21x2_ASAP7_75t_L g677 ( .A1(n_634), .A2(n_151), .B(n_235), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_540), .Y(n_678) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_626), .A2(n_150), .B(n_234), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_583), .Y(n_680) );
OA21x2_ASAP7_75t_L g681 ( .A1(n_593), .A2(n_148), .B(n_233), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_555), .B(n_34), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_535), .B(n_35), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_603), .A2(n_145), .B(n_228), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_612), .A2(n_144), .B(n_227), .Y(n_685) );
OAI22xp33_ASAP7_75t_SL g686 ( .A1(n_564), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_686) );
OAI21x1_ASAP7_75t_L g687 ( .A1(n_570), .A2(n_157), .B(n_226), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_623), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_627), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_640), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_572), .B(n_38), .Y(n_691) );
CKINVDCx8_ASAP7_75t_R g692 ( .A(n_580), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_547), .B(n_38), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_549), .Y(n_694) );
OAI21x1_ASAP7_75t_L g695 ( .A1(n_582), .A2(n_142), .B(n_222), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_608), .B(n_40), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_632), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_578), .A2(n_41), .B(n_42), .C(n_43), .Y(n_698) );
OA21x2_ASAP7_75t_L g699 ( .A1(n_575), .A2(n_159), .B(n_221), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_582), .A2(n_141), .B(n_220), .Y(n_700) );
OAI21x1_ASAP7_75t_L g701 ( .A1(n_638), .A2(n_139), .B(n_219), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_539), .B(n_42), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_641), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_584), .Y(n_704) );
OAI21x1_ASAP7_75t_L g705 ( .A1(n_551), .A2(n_160), .B(n_218), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_619), .A2(n_135), .B(n_216), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_587), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_563), .Y(n_708) );
BUFx3_ASAP7_75t_L g709 ( .A(n_599), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_L g710 ( .A1(n_573), .A2(n_43), .B(n_44), .C(n_45), .Y(n_710) );
INVx4_ASAP7_75t_L g711 ( .A(n_618), .Y(n_711) );
NAND2xp33_ASAP7_75t_L g712 ( .A(n_632), .B(n_590), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_532), .B(n_47), .Y(n_713) );
OA21x2_ASAP7_75t_L g714 ( .A1(n_629), .A2(n_164), .B(n_211), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_635), .A2(n_47), .B1(n_49), .B2(n_50), .Y(n_715) );
OA21x2_ASAP7_75t_L g716 ( .A1(n_562), .A2(n_168), .B(n_210), .Y(n_716) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_565), .A2(n_161), .B(n_207), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_624), .Y(n_718) );
AO21x2_ASAP7_75t_L g719 ( .A1(n_615), .A2(n_134), .B(n_206), .Y(n_719) );
OA21x2_ASAP7_75t_L g720 ( .A1(n_628), .A2(n_129), .B(n_204), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_571), .A2(n_50), .B1(n_51), .B2(n_53), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_588), .A2(n_51), .B1(n_53), .B2(n_55), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_563), .Y(n_723) );
OA21x2_ASAP7_75t_L g724 ( .A1(n_561), .A2(n_170), .B(n_201), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_563), .Y(n_725) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_635), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_577), .A2(n_56), .B(n_57), .C(n_58), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_611), .A2(n_116), .B(n_199), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_542), .B(n_56), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_548), .B(n_57), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_614), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_602), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_633), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_553), .B(n_58), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_548), .B(n_59), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_552), .B(n_60), .Y(n_736) );
NOR2x1_ASAP7_75t_R g737 ( .A(n_553), .B(n_62), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_594), .Y(n_738) );
OAI21x1_ASAP7_75t_L g739 ( .A1(n_569), .A2(n_96), .B(n_97), .Y(n_739) );
AO21x2_ASAP7_75t_L g740 ( .A1(n_585), .A2(n_101), .B(n_105), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_541), .A2(n_108), .B1(n_109), .B2(n_113), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_589), .Y(n_742) );
AO31x2_ASAP7_75t_L g743 ( .A1(n_625), .A2(n_242), .A3(n_176), .B(n_178), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_585), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_589), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_560), .Y(n_746) );
INVx2_ASAP7_75t_SL g747 ( .A(n_620), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_557), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_595), .A2(n_173), .B1(n_180), .B2(n_182), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_595), .A2(n_183), .B1(n_187), .B2(n_188), .Y(n_750) );
BUFx4f_ASAP7_75t_SL g751 ( .A(n_694), .Y(n_751) );
NOR4xp25_ASAP7_75t_L g752 ( .A(n_668), .B(n_621), .C(n_537), .D(n_597), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_646), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_744), .A2(n_607), .B1(n_554), .B2(n_574), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_703), .A2(n_591), .B(n_605), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_696), .A2(n_609), .B1(n_543), .B2(n_591), .C(n_531), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_704), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_744), .A2(n_545), .B1(n_536), .B2(n_544), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_712), .A2(n_637), .B(n_631), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_670), .B(n_682), .Y(n_760) );
INVx3_ASAP7_75t_L g761 ( .A(n_711), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_712), .A2(n_637), .B(n_631), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_668), .A2(n_598), .B1(n_590), .B2(n_568), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_658), .A2(n_728), .B(n_684), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_651), .B(n_191), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_696), .B(n_196), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_689), .A2(n_198), .B1(n_726), .B2(n_676), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_662), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_659), .A2(n_736), .B1(n_730), .B2(n_735), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_693), .B(n_683), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_661), .B(n_738), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_676), .B(n_654), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_704), .A2(n_736), .B1(n_729), .B2(n_707), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_721), .A2(n_731), .B(n_671), .Y(n_774) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_691), .A2(n_702), .B(n_678), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_663), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_673), .B(n_713), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_662), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_650), .B(n_690), .Y(n_779) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_710), .A2(n_747), .B1(n_749), .B2(n_750), .C(n_653), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_708), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_749), .A2(n_750), .B1(n_715), .B2(n_669), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_655), .A2(n_665), .B(n_675), .Y(n_783) );
OA21x2_ASAP7_75t_L g784 ( .A1(n_655), .A2(n_657), .B(n_706), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_694), .Y(n_785) );
AOI211xp5_ASAP7_75t_L g786 ( .A1(n_737), .A2(n_686), .B(n_734), .C(n_727), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_643), .A2(n_647), .B1(n_667), .B2(n_722), .Y(n_787) );
AO221x2_ASAP7_75t_L g788 ( .A1(n_666), .A2(n_742), .B1(n_745), .B2(n_644), .C(n_698), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_649), .B(n_732), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_665), .A2(n_675), .B(n_714), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_709), .B(n_656), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_746), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_748), .Y(n_793) );
OAI221xp5_ASAP7_75t_SL g794 ( .A1(n_645), .A2(n_741), .B1(n_725), .B2(n_723), .C(n_708), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_680), .B(n_723), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_718), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_652), .B(n_725), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_644), .B(n_652), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_733), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_644), .B(n_652), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_646), .B(n_688), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_665), .A2(n_675), .B(n_714), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_740), .A2(n_720), .B1(n_724), .B2(n_681), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_743), .B(n_688), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_743), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_701), .A2(n_685), .B(n_687), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_720), .A2(n_724), .B1(n_681), .B2(n_719), .Y(n_807) );
AO221x2_ASAP7_75t_L g808 ( .A1(n_743), .A2(n_692), .B1(n_681), .B2(n_714), .C(n_664), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_672), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_677), .A2(n_699), .B(n_717), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_646), .A2(n_724), .B1(n_697), .B2(n_672), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_674), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_660), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_664), .A2(n_699), .B1(n_716), .B2(n_717), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_743), .Y(n_815) );
OAI221xp5_ASAP7_75t_L g816 ( .A1(n_705), .A2(n_679), .B1(n_648), .B2(n_739), .C(n_695), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_679), .B(n_700), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_642), .A2(n_744), .B1(n_571), .B2(n_668), .Y(n_818) );
NAND2x1_ASAP7_75t_L g819 ( .A(n_711), .B(n_583), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_651), .B(n_448), .Y(n_820) );
OR2x6_ASAP7_75t_L g821 ( .A(n_676), .B(n_540), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_703), .A2(n_630), .B(n_558), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_711), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_704), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_651), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_651), .B(n_448), .Y(n_826) );
BUFx2_ASAP7_75t_L g827 ( .A(n_704), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_744), .A2(n_571), .B1(n_555), .B2(n_576), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_704), .Y(n_829) );
CKINVDCx11_ASAP7_75t_R g830 ( .A(n_692), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_651), .B(n_448), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_662), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_670), .B(n_448), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_744), .A2(n_454), .B1(n_670), .B2(n_571), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_651), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_662), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_651), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_744), .A2(n_689), .B1(n_726), .B2(n_433), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_744), .A2(n_571), .B1(n_555), .B2(n_576), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_744), .B(n_639), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_768), .B(n_778), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_832), .B(n_836), .Y(n_842) );
INVxp67_ASAP7_75t_L g843 ( .A(n_757), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_797), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_804), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_821), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_813), .Y(n_847) );
INVx3_ASAP7_75t_L g848 ( .A(n_753), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_798), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_800), .Y(n_850) );
AO21x2_ASAP7_75t_L g851 ( .A1(n_790), .A2(n_802), .B(n_783), .Y(n_851) );
OR2x2_ASAP7_75t_L g852 ( .A(n_769), .B(n_770), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_776), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_833), .B(n_760), .Y(n_854) );
BUFx3_ASAP7_75t_L g855 ( .A(n_819), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_825), .B(n_835), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_837), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_796), .B(n_799), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_793), .B(n_792), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_769), .B(n_781), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_838), .B(n_840), .Y(n_861) );
AND2x4_ASAP7_75t_SL g862 ( .A(n_761), .B(n_823), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_805), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_815), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_817), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_834), .A2(n_786), .B1(n_773), .B2(n_782), .C(n_752), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_820), .B(n_826), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_777), .B(n_791), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_751), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_828), .B(n_839), .Y(n_870) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_775), .A2(n_767), .B(n_772), .C(n_794), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_788), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_831), .B(n_771), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_795), .B(n_788), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_812), .B(n_766), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_818), .B(n_774), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_751), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_784), .Y(n_878) );
BUFx2_ASAP7_75t_L g879 ( .A(n_801), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_808), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_809), .B(n_806), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_789), .Y(n_882) );
NOR4xp25_ASAP7_75t_SL g883 ( .A(n_780), .B(n_816), .C(n_827), .D(n_824), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_754), .A2(n_787), .B1(n_763), .B2(n_756), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_779), .B(n_763), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_755), .B(n_765), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_808), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_784), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_758), .B(n_759), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_759), .B(n_762), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_785), .A2(n_829), .B1(n_764), .B2(n_830), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_803), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_807), .B(n_762), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_811), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_807), .B(n_814), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_814), .Y(n_896) );
INVx4_ASAP7_75t_L g897 ( .A(n_822), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_802), .B(n_810), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_863), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_849), .B(n_850), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_864), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_868), .B(n_850), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_895), .B(n_872), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_872), .B(n_874), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_874), .B(n_896), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_896), .B(n_865), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_860), .B(n_844), .Y(n_907) );
OAI211xp5_ASAP7_75t_SL g908 ( .A1(n_843), .A2(n_891), .B(n_866), .C(n_867), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_841), .B(n_842), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_841), .B(n_842), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_854), .B(n_880), .Y(n_911) );
OAI322xp33_ASAP7_75t_L g912 ( .A1(n_860), .A2(n_891), .A3(n_861), .B1(n_852), .B2(n_870), .C1(n_873), .C2(n_884), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_887), .B(n_856), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_887), .B(n_856), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_852), .B(n_870), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_845), .B(n_859), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_871), .A2(n_846), .B1(n_882), .B2(n_857), .C(n_853), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_875), .A2(n_885), .B1(n_876), .B2(n_882), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_859), .B(n_858), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_892), .B(n_893), .Y(n_920) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_869), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_858), .B(n_892), .Y(n_922) );
OAI221xp5_ASAP7_75t_SL g923 ( .A1(n_889), .A2(n_893), .B1(n_877), .B2(n_875), .C(n_890), .Y(n_923) );
INVx4_ASAP7_75t_L g924 ( .A(n_855), .Y(n_924) );
INVx3_ASAP7_75t_L g925 ( .A(n_881), .Y(n_925) );
INVx4_ASAP7_75t_L g926 ( .A(n_855), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_886), .B(n_879), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_921), .B(n_862), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_919), .B(n_862), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_905), .B(n_881), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_899), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_899), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_906), .B(n_851), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_901), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_906), .B(n_851), .Y(n_935) );
NOR3xp33_ASAP7_75t_SL g936 ( .A(n_908), .B(n_883), .C(n_897), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_903), .B(n_847), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_927), .B(n_898), .Y(n_938) );
INVx3_ASAP7_75t_L g939 ( .A(n_924), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_927), .B(n_894), .Y(n_940) );
NOR2xp67_ASAP7_75t_SL g941 ( .A(n_917), .B(n_848), .Y(n_941) );
BUFx2_ASAP7_75t_L g942 ( .A(n_924), .Y(n_942) );
INVx1_ASAP7_75t_SL g943 ( .A(n_909), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_900), .B(n_878), .Y(n_944) );
AND2x4_ASAP7_75t_L g945 ( .A(n_925), .B(n_897), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_900), .B(n_878), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_904), .B(n_888), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_904), .B(n_888), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_943), .B(n_907), .Y(n_949) );
AOI211xp5_ASAP7_75t_L g950 ( .A1(n_941), .A2(n_912), .B(n_923), .C(n_918), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_933), .B(n_925), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_935), .B(n_925), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_931), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_935), .B(n_920), .Y(n_954) );
OR2x6_ASAP7_75t_L g955 ( .A(n_942), .B(n_926), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_932), .Y(n_956) );
INVx1_ASAP7_75t_SL g957 ( .A(n_929), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_940), .B(n_920), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_928), .B(n_911), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_932), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_940), .B(n_915), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_934), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_939), .Y(n_963) );
INVx3_ASAP7_75t_SL g964 ( .A(n_939), .Y(n_964) );
NAND2x1p5_ASAP7_75t_L g965 ( .A(n_963), .B(n_926), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g966 ( .A1(n_963), .A2(n_918), .B1(n_939), .B2(n_911), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g967 ( .A(n_950), .B(n_941), .C(n_936), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_949), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_949), .B(n_938), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_959), .A2(n_913), .B1(n_914), .B2(n_902), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_969), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_966), .A2(n_964), .B1(n_955), .B2(n_961), .Y(n_972) );
XNOR2xp5_ASAP7_75t_L g973 ( .A(n_967), .B(n_957), .Y(n_973) );
OAI22xp33_ASAP7_75t_SL g974 ( .A1(n_965), .A2(n_955), .B1(n_958), .B2(n_926), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_968), .B(n_954), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_972), .A2(n_970), .B1(n_952), .B2(n_951), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_975), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_973), .A2(n_930), .B1(n_947), .B2(n_948), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_974), .A2(n_944), .B(n_946), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_971), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_976), .A2(n_978), .B1(n_977), .B2(n_980), .Y(n_981) );
AOI321xp33_ASAP7_75t_L g982 ( .A1(n_979), .A2(n_937), .A3(n_945), .B1(n_962), .B2(n_960), .C(n_956), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_981), .B(n_962), .Y(n_983) );
INVx4_ASAP7_75t_L g984 ( .A(n_982), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_983), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_984), .B(n_953), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_986), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_985), .Y(n_988) );
INVx4_ASAP7_75t_L g989 ( .A(n_988), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_987), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_989), .Y(n_991) );
NAND2xp33_ASAP7_75t_SL g992 ( .A(n_991), .B(n_990), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_992), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_993), .A2(n_922), .B1(n_910), .B2(n_916), .Y(n_994) );
endmodule