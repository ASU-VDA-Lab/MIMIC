module fake_jpeg_6529_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_37),
.B(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_38),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_0),
.B(n_2),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_28),
.C(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_21),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_24),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_54),
.B(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_64),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_71),
.B1(n_85),
.B2(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_70),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_25),
.B1(n_35),
.B2(n_18),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_93),
.B1(n_19),
.B2(n_34),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_30),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_77),
.Y(n_119)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_74),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_84),
.Y(n_111)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_39),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_40),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_22),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_21),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_74),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_20),
.B1(n_19),
.B2(n_21),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_121),
.B1(n_124),
.B2(n_6),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_76),
.B1(n_116),
.B2(n_8),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_85),
.B1(n_62),
.B2(n_71),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_147),
.B1(n_109),
.B2(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_98),
.B1(n_81),
.B2(n_83),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_125),
.B1(n_109),
.B2(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_55),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_143),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_53),
.C(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_70),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_81),
.B1(n_79),
.B2(n_76),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_60),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_156),
.B1(n_116),
.B2(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_157),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_94),
.B(n_96),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_158),
.B(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_99),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_7),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_7),
.B(n_8),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_172),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_112),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_83),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_183),
.B1(n_184),
.B2(n_129),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_137),
.B1(n_134),
.B2(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_101),
.C(n_113),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_157),
.C(n_158),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_123),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_178),
.B(n_11),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_101),
.B(n_103),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_127),
.B1(n_108),
.B2(n_113),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_108),
.B1(n_105),
.B2(n_103),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_105),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_155),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_198),
.B(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_205),
.C(n_206),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_203),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_161),
.B1(n_180),
.B2(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_186),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_8),
.B(n_9),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_140),
.B(n_146),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_11),
.C(n_12),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_11),
.C(n_160),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_219),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_173),
.B1(n_167),
.B2(n_165),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_201),
.B1(n_188),
.B2(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_188),
.B1(n_197),
.B2(n_165),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_202),
.B1(n_169),
.B2(n_168),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_175),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_215),
.B1(n_184),
.B2(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_219),
.C(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_233),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_201),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_211),
.C(n_210),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_211),
.C(n_190),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_179),
.C(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_245),
.B(n_166),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_226),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_248),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

AOI31xp33_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_218),
.A3(n_207),
.B(n_216),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_230),
.A3(n_231),
.B1(n_229),
.B2(n_198),
.C1(n_159),
.C2(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_163),
.B(n_200),
.Y(n_263)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_181),
.B(n_204),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_215),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_234),
.B1(n_204),
.B2(n_164),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_247),
.B(n_250),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_259),
.B(n_253),
.C(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_256),
.B(n_254),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_266),
.B(n_159),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_205),
.CI(n_178),
.CON(n_267),
.SN(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_268),
.Y(n_270)
);


endmodule