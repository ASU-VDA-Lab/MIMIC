module real_aes_16696_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g112 ( .A(n_0), .B(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_1), .A2(n_4), .B1(n_277), .B2(n_278), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_2), .A2(n_43), .B1(n_178), .B2(n_226), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_3), .A2(n_24), .B1(n_226), .B2(n_260), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_5), .A2(n_16), .B1(n_527), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_6), .A2(n_62), .B1(n_163), .B2(n_164), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_7), .A2(n_17), .B1(n_178), .B2(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_9), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_10), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_11), .A2(n_18), .B1(n_528), .B2(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_12), .A2(n_66), .B1(n_136), .B2(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
OR2x2_ASAP7_75t_L g108 ( .A(n_13), .B(n_38), .Y(n_108) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_15), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_19), .A2(n_99), .B1(n_278), .B2(n_527), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_20), .A2(n_39), .B1(n_156), .B2(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_21), .B(n_154), .Y(n_588) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_22), .A2(n_59), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_23), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_25), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_26), .B(n_151), .Y(n_218) );
INVx4_ASAP7_75t_R g202 ( .A(n_27), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_28), .A2(n_47), .B1(n_182), .B2(n_275), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_29), .A2(n_54), .B1(n_182), .B2(n_527), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_30), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_31), .B(n_552), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_32), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_33), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g282 ( .A(n_34), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_SL g257 ( .A1(n_35), .A2(n_150), .B(n_178), .C(n_258), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_36), .A2(n_55), .B1(n_178), .B2(n_182), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_37), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_40), .A2(n_87), .B1(n_178), .B2(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g822 ( .A1(n_41), .A2(n_53), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_41), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_42), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_44), .A2(n_46), .B1(n_178), .B2(n_179), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_45), .A2(n_60), .B1(n_527), .B2(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g222 ( .A(n_48), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_49), .B(n_178), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_50), .Y(n_236) );
INVx2_ASAP7_75t_L g131 ( .A(n_51), .Y(n_131) );
BUFx3_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
INVx1_ASAP7_75t_L g125 ( .A(n_52), .Y(n_125) );
INVx1_ASAP7_75t_L g823 ( .A(n_53), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_56), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_57), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_58), .A2(n_88), .B1(n_178), .B2(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g826 ( .A(n_61), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_63), .A2(n_76), .B1(n_275), .B2(n_544), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_64), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_65), .A2(n_79), .B1(n_178), .B2(n_179), .Y(n_529) );
INVx1_ASAP7_75t_L g137 ( .A(n_66), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_67), .A2(n_98), .B1(n_527), .B2(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g169 ( .A(n_68), .Y(n_169) );
AND2x4_ASAP7_75t_L g172 ( .A(n_69), .B(n_173), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_70), .A2(n_90), .B1(n_182), .B2(n_275), .Y(n_274) );
AO22x1_ASAP7_75t_L g152 ( .A1(n_71), .A2(n_77), .B1(n_153), .B2(n_156), .Y(n_152) );
INVx1_ASAP7_75t_L g173 ( .A(n_72), .Y(n_173) );
AND2x2_ASAP7_75t_L g261 ( .A(n_73), .B(n_214), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_74), .B(n_163), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_75), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_78), .B(n_226), .Y(n_237) );
INVx2_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_81), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_82), .B(n_214), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_83), .A2(n_97), .B1(n_163), .B2(n_182), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_84), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_85), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_86), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_89), .B(n_214), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_91), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_92), .B(n_214), .Y(n_233) );
INVx1_ASAP7_75t_L g111 ( .A(n_93), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_93), .B(n_124), .Y(n_123) );
NAND2xp33_ASAP7_75t_L g591 ( .A(n_94), .B(n_154), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_95), .A2(n_163), .B(n_184), .C(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g207 ( .A(n_96), .B(n_208), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g241 ( .A(n_100), .B(n_203), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_114), .B(n_825), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
BUFx12f_ASAP7_75t_L g828 ( .A(n_104), .Y(n_828) );
OR2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_109), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g810 ( .A(n_106), .B(n_499), .Y(n_810) );
NOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g133 ( .A(n_107), .Y(n_133) );
INVx1_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g499 ( .A(n_111), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g114 ( .A(n_115), .B(n_811), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_127), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_117), .A2(n_817), .B(n_819), .Y(n_816) );
NOR2x1_ASAP7_75t_R g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g818 ( .A(n_120), .Y(n_818) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_126), .B(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_804), .Y(n_127) );
BUFx12f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x6_ASAP7_75t_SL g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_131), .B(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g815 ( .A(n_131), .Y(n_815) );
OAI22xp33_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_138), .B1(n_139), .B2(n_803), .Y(n_134) );
INVx1_ASAP7_75t_L g803 ( .A(n_135), .Y(n_803) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_497), .B1(n_500), .B2(n_802), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_407), .Y(n_141) );
NOR3xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_336), .C(n_378), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_310), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_209), .B1(n_285), .B2(n_296), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_190), .Y(n_146) );
AOI21xp33_ASAP7_75t_L g329 ( .A1(n_147), .A2(n_330), .B(n_332), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_147), .A2(n_403), .B(n_404), .Y(n_402) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_174), .Y(n_147) );
INVx2_ASAP7_75t_L g322 ( .A(n_148), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_148), .B(n_175), .Y(n_352) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_158), .C(n_170), .Y(n_149) );
INVx6_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_150), .A2(n_241), .B(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_150), .B(n_152), .Y(n_294) );
O2A1O1Ixp5_ASAP7_75t_L g586 ( .A1(n_150), .A2(n_179), .B(n_587), .C(n_588), .Y(n_586) );
BUFx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
INVx1_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
INVxp67_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g527 ( .A(n_154), .Y(n_527) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g157 ( .A(n_155), .Y(n_157) );
INVx1_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_155), .Y(n_165) );
INVx3_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g254 ( .A(n_155), .Y(n_254) );
INVx2_ASAP7_75t_L g260 ( .A(n_155), .Y(n_260) );
OAI21xp33_ASAP7_75t_SL g217 ( .A1(n_156), .A2(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g293 ( .A(n_158), .Y(n_293) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_166), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_159), .A2(n_224), .B(n_225), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_159), .A2(n_180), .B1(n_265), .B2(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g510 ( .A(n_160), .Y(n_510) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
INVx1_ASAP7_75t_L g572 ( .A(n_164), .Y(n_572) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_199), .Y(n_198) );
OAI21xp33_ASAP7_75t_L g170 ( .A1(n_166), .A2(n_167), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVx2_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
INVx1_ASAP7_75t_L g295 ( .A(n_170), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_171), .A2(n_250), .B(n_257), .Y(n_249) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx10_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
BUFx10_ASAP7_75t_L g228 ( .A(n_172), .Y(n_228) );
INVx1_ASAP7_75t_L g280 ( .A(n_172), .Y(n_280) );
AND2x2_ASAP7_75t_L g392 ( .A(n_174), .B(n_231), .Y(n_392) );
INVx1_ASAP7_75t_L g425 ( .A(n_174), .Y(n_425) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g287 ( .A(n_175), .B(n_232), .Y(n_287) );
AND2x2_ASAP7_75t_L g318 ( .A(n_175), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g327 ( .A(n_175), .Y(n_327) );
OR2x2_ASAP7_75t_L g346 ( .A(n_175), .B(n_192), .Y(n_346) );
AND2x2_ASAP7_75t_L g361 ( .A(n_175), .B(n_192), .Y(n_361) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_185), .A3(n_186), .B(n_187), .Y(n_175) );
OAI22x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B1(n_181), .B2(n_183), .Y(n_176) );
INVx4_ASAP7_75t_L g179 ( .A(n_178), .Y(n_179) );
INVx1_ASAP7_75t_L g528 ( .A(n_178), .Y(n_528) );
INVx1_ASAP7_75t_L g544 ( .A(n_178), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_179), .A2(n_236), .B(n_237), .C(n_238), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_180), .A2(n_183), .B1(n_274), .B2(n_276), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_180), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_180), .A2(n_183), .B1(n_518), .B2(n_520), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_180), .A2(n_526), .B1(n_529), .B2(n_530), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_180), .A2(n_510), .B1(n_542), .B2(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_180), .A2(n_510), .B1(n_551), .B2(n_553), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_180), .A2(n_510), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_180), .A2(n_530), .B1(n_571), .B2(n_573), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_180), .A2(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_182), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g277 ( .A(n_182), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_183), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_SL g530 ( .A(n_184), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_185), .B(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_185), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g206 ( .A(n_186), .Y(n_206) );
AO31x2_ASAP7_75t_L g507 ( .A1(n_186), .A2(n_267), .A3(n_508), .B(n_512), .Y(n_507) );
AO31x2_ASAP7_75t_L g549 ( .A1(n_186), .A2(n_516), .A3(n_550), .B(n_555), .Y(n_549) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_186), .A2(n_248), .A3(n_570), .B(n_574), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx2_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
BUFx2_ASAP7_75t_L g248 ( .A(n_189), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_189), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_189), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_191), .B(n_360), .Y(n_403) );
OR2x2_ASAP7_75t_L g491 ( .A(n_191), .B(n_352), .Y(n_491) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g319 ( .A(n_192), .Y(n_319) );
AND2x2_ASAP7_75t_L g328 ( .A(n_192), .B(n_291), .Y(n_328) );
AND2x2_ASAP7_75t_L g331 ( .A(n_192), .B(n_232), .Y(n_331) );
AND2x2_ASAP7_75t_L g350 ( .A(n_192), .B(n_231), .Y(n_350) );
AND2x4_ASAP7_75t_L g369 ( .A(n_192), .B(n_292), .Y(n_369) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_196), .B(n_207), .Y(n_192) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_193), .A2(n_531), .A3(n_541), .B(n_545), .Y(n_540) );
AO31x2_ASAP7_75t_L g559 ( .A1(n_193), .A2(n_279), .A3(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_195), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_SL g574 ( .A(n_195), .B(n_575), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_200), .B(n_206), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_201) );
INVx2_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
INVx1_ASAP7_75t_L g552 ( .A(n_203), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_204), .Y(n_554) );
INVx1_ASAP7_75t_L g531 ( .A(n_206), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_229), .B(n_270), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_210), .B(n_364), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_212), .B(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g300 ( .A(n_212), .Y(n_300) );
OR2x2_ASAP7_75t_L g308 ( .A(n_212), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_212), .B(n_301), .Y(n_333) );
AND2x2_ASAP7_75t_L g358 ( .A(n_212), .B(n_272), .Y(n_358) );
AND2x2_ASAP7_75t_L g376 ( .A(n_212), .B(n_306), .Y(n_376) );
INVx1_ASAP7_75t_L g415 ( .A(n_212), .Y(n_415) );
AND2x2_ASAP7_75t_L g417 ( .A(n_212), .B(n_418), .Y(n_417) );
NAND2x1p5_ASAP7_75t_SL g436 ( .A(n_212), .B(n_357), .Y(n_436) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_216), .Y(n_212) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_214), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g227 ( .A(n_215), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_215), .B(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g516 ( .A(n_215), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_215), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_215), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g584 ( .A(n_215), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_223), .B(n_227), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
BUFx4f_ASAP7_75t_L g256 ( .A(n_221), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_226), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_228), .A2(n_264), .A3(n_267), .B(n_268), .Y(n_263) );
OAI32xp33_ASAP7_75t_L g320 ( .A1(n_229), .A2(n_312), .A3(n_321), .B1(n_323), .B2(n_325), .Y(n_320) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_245), .Y(n_229) );
INVx1_ASAP7_75t_L g360 ( .A(n_230), .Y(n_360) );
AND2x2_ASAP7_75t_L g368 ( .A(n_230), .B(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g367 ( .A(n_231), .B(n_291), .Y(n_367) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
BUFx3_ASAP7_75t_L g317 ( .A(n_232), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g432 ( .A(n_232), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_240), .B(n_243), .Y(n_234) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g302 ( .A(n_245), .Y(n_302) );
OR2x2_ASAP7_75t_L g312 ( .A(n_245), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g434 ( .A(n_245), .Y(n_434) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_262), .Y(n_245) );
AND2x2_ASAP7_75t_L g335 ( .A(n_246), .B(n_263), .Y(n_335) );
INVx2_ASAP7_75t_L g357 ( .A(n_246), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_246), .B(n_272), .Y(n_377) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g284 ( .A(n_247), .Y(n_284) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_261), .Y(n_247) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_248), .A2(n_273), .A3(n_279), .B(n_281), .Y(n_272) );
AO31x2_ASAP7_75t_L g524 ( .A1(n_248), .A2(n_525), .A3(n_531), .B(n_532), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B(n_256), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_SL g519 ( .A(n_260), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_262), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g366 ( .A(n_262), .Y(n_366) );
INVx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
OR2x2_ASAP7_75t_L g372 ( .A(n_263), .B(n_272), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_263), .B(n_272), .Y(n_405) );
INVx2_ASAP7_75t_L g353 ( .A(n_270), .Y(n_353) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_283), .Y(n_270) );
OR2x2_ASAP7_75t_L g340 ( .A(n_271), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g418 ( .A(n_271), .Y(n_418) );
INVx1_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
INVx1_ASAP7_75t_L g309 ( .A(n_272), .Y(n_309) );
INVx1_ASAP7_75t_L g324 ( .A(n_272), .Y(n_324) );
AO31x2_ASAP7_75t_L g515 ( .A1(n_279), .A2(n_516), .A3(n_517), .B(n_521), .Y(n_515) );
INVx2_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g592 ( .A(n_280), .Y(n_592) );
OR2x2_ASAP7_75t_L g428 ( .A(n_283), .B(n_405), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_284), .B(n_300), .Y(n_341) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_284), .Y(n_343) );
OR2x2_ASAP7_75t_L g442 ( .A(n_284), .B(n_366), .Y(n_442) );
INVxp67_ASAP7_75t_L g466 ( .A(n_284), .Y(n_466) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_287), .B(n_328), .Y(n_395) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g344 ( .A(n_289), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g457 ( .A(n_290), .Y(n_457) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g486 ( .A(n_291), .B(n_319), .Y(n_486) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g412 ( .A(n_292), .B(n_319), .Y(n_412) );
AOI21x1_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_303), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_299), .B(n_335), .Y(n_449) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
AND2x2_ASAP7_75t_L g363 ( .A(n_300), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_300), .B(n_357), .Y(n_406) );
OR2x2_ASAP7_75t_L g478 ( .A(n_300), .B(n_365), .Y(n_478) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_304), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx2_ASAP7_75t_L g389 ( .A(n_305), .Y(n_389) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g379 ( .A(n_308), .B(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_308), .Y(n_390) );
OR2x2_ASAP7_75t_L g441 ( .A(n_308), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g496 ( .A(n_308), .Y(n_496) );
AOI211xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_320), .C(n_329), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g385 ( .A(n_313), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_313), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g458 ( .A(n_313), .B(n_335), .Y(n_458) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_316), .B(n_361), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_316), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g468 ( .A(n_316), .B(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g411 ( .A(n_317), .Y(n_411) );
AND2x2_ASAP7_75t_L g439 ( .A(n_318), .B(n_367), .Y(n_439) );
INVx2_ASAP7_75t_L g462 ( .A(n_318), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_318), .B(n_360), .Y(n_494) );
AND2x4_ASAP7_75t_SL g448 ( .A(n_321), .B(n_326), .Y(n_448) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g401 ( .A(n_322), .B(n_327), .Y(n_401) );
OR2x2_ASAP7_75t_L g453 ( .A(n_322), .B(n_346), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_323), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_323), .B(n_335), .Y(n_489) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g437 ( .A(n_324), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g420 ( .A(n_326), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_326), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g470 ( .A(n_327), .Y(n_470) );
BUFx2_ASAP7_75t_L g338 ( .A(n_328), .Y(n_338) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g456 ( .A(n_331), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_335), .Y(n_397) );
NAND3xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_347), .C(n_362), .Y(n_336) );
AOI22xp33_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_339), .B1(n_342), .B2(n_344), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_344), .A2(n_370), .B1(n_451), .B2(n_454), .C1(n_456), .C2(n_458), .Y(n_450) );
AND2x2_ASAP7_75t_L g482 ( .A(n_345), .B(n_431), .Y(n_482) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g430 ( .A(n_346), .B(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_353), .B1(n_354), .B2(n_359), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_SL g426 ( .A(n_350), .Y(n_426) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
AND2x2_ASAP7_75t_L g413 ( .A(n_355), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g371 ( .A(n_356), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g365 ( .A(n_357), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g480 ( .A(n_358), .Y(n_480) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_361), .B(n_457), .Y(n_476) );
INVx1_ASAP7_75t_L g493 ( .A(n_361), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_368), .B2(n_370), .C1(n_373), .C2(n_374), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_369), .Y(n_373) );
AND2x2_ASAP7_75t_L g391 ( .A(n_369), .B(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g422 ( .A(n_369), .Y(n_422) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g386 ( .A(n_372), .Y(n_386) );
OR2x2_ASAP7_75t_L g455 ( .A(n_372), .B(n_436), .Y(n_455) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_384), .C(n_393), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_391), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_385), .A2(n_423), .B1(n_472), .B2(n_475), .C(n_477), .Y(n_471) );
AND2x4_ASAP7_75t_L g414 ( .A(n_386), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
AOI211x1_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_398), .C(n_402), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g463 ( .A(n_401), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_404), .B(n_452), .C(n_453), .Y(n_451) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_459), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_416), .C(n_438), .D(n_450), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
AND2x2_ASAP7_75t_L g469 ( .A(n_412), .B(n_470), .Y(n_469) );
AOI221x1_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_439), .B1(n_440), .B2(n_443), .C(n_446), .Y(n_438) );
AND2x2_ASAP7_75t_L g464 ( .A(n_414), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g474 ( .A(n_415), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_423), .B2(n_427), .C(n_429), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_421), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_426), .A2(n_430), .B1(n_433), .B2(n_435), .Y(n_429) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_430), .A2(n_447), .B(n_449), .Y(n_446) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g473 ( .A(n_442), .Y(n_473) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_455), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_483), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B1(n_467), .B2(n_468), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g479 ( .A(n_466), .B(n_480), .Y(n_479) );
NAND2x1_ASAP7_75t_L g495 ( .A(n_466), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_481), .Y(n_477) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B1(n_488), .B2(n_490), .C(n_492), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g802 ( .A(n_497), .Y(n_802) );
BUFx12f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_500), .B(n_822), .Y(n_821) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_501), .B(n_712), .Y(n_500) );
NAND4xp75_ASAP7_75t_L g501 ( .A(n_502), .B(n_657), .C(n_677), .D(n_693), .Y(n_501) );
NOR2x1p5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_627), .Y(n_502) );
NAND4xp75_ASAP7_75t_L g503 ( .A(n_504), .B(n_565), .C(n_604), .D(n_613), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_534), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
AND2x4_ASAP7_75t_L g737 ( .A(n_506), .B(n_664), .Y(n_737) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_507), .Y(n_580) );
INVx2_ASAP7_75t_L g598 ( .A(n_507), .Y(n_598) );
AND2x2_ASAP7_75t_L g621 ( .A(n_507), .B(n_583), .Y(n_621) );
OR2x2_ASAP7_75t_L g676 ( .A(n_507), .B(n_515), .Y(n_676) );
AND2x2_ASAP7_75t_L g594 ( .A(n_514), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g744 ( .A(n_514), .B(n_621), .Y(n_744) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
OR2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g612 ( .A(n_515), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_515), .B(n_524), .Y(n_618) );
INVx1_ASAP7_75t_L g636 ( .A(n_515), .Y(n_636) );
INVx2_ASAP7_75t_L g665 ( .A(n_515), .Y(n_665) );
INVx3_ASAP7_75t_L g641 ( .A(n_523), .Y(n_641) );
INVx2_ASAP7_75t_L g646 ( .A(n_523), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_523), .B(n_597), .Y(n_651) );
AND2x2_ASAP7_75t_L g674 ( .A(n_523), .B(n_653), .Y(n_674) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_523), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_523), .B(n_729), .Y(n_728) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g663 ( .A(n_524), .Y(n_663) );
AND2x2_ASAP7_75t_L g711 ( .A(n_524), .B(n_665), .Y(n_711) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_547), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_536), .B(n_655), .Y(n_702) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g699 ( .A(n_537), .B(n_655), .Y(n_699) );
INVx1_ASAP7_75t_L g800 ( .A(n_537), .Y(n_800) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g750 ( .A(n_538), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
OR2x2_ASAP7_75t_L g684 ( .A(n_539), .B(n_558), .Y(n_684) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g626 ( .A(n_540), .Y(n_626) );
AND2x4_ASAP7_75t_L g632 ( .A(n_540), .B(n_633), .Y(n_632) );
AOI32xp33_ASAP7_75t_L g770 ( .A1(n_547), .A2(n_673), .A3(n_771), .B1(n_773), .B2(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g719 ( .A(n_548), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_557), .Y(n_548) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_549), .Y(n_567) );
OR2x2_ASAP7_75t_L g601 ( .A(n_549), .B(n_559), .Y(n_601) );
INVx1_ASAP7_75t_L g616 ( .A(n_549), .Y(n_616) );
AND2x2_ASAP7_75t_L g625 ( .A(n_549), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g631 ( .A(n_549), .Y(n_631) );
INVx2_ASAP7_75t_L g656 ( .A(n_549), .Y(n_656) );
AND2x2_ASAP7_75t_L g775 ( .A(n_549), .B(n_569), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_557), .B(n_608), .Y(n_695) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g568 ( .A(n_559), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g624 ( .A(n_559), .Y(n_624) );
INVx2_ASAP7_75t_L g633 ( .A(n_559), .Y(n_633) );
AND2x4_ASAP7_75t_L g655 ( .A(n_559), .B(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_559), .Y(n_747) );
AOI22x1_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_576), .B1(n_594), .B2(n_599), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_568), .B(n_725), .C(n_726), .D(n_727), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_568), .B(n_625), .Y(n_755) );
INVx4_ASAP7_75t_SL g608 ( .A(n_569), .Y(n_608) );
BUFx2_ASAP7_75t_L g671 ( .A(n_569), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_569), .B(n_616), .Y(n_734) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g696 ( .A(n_578), .B(n_645), .Y(n_696) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g619 ( .A(n_582), .B(n_597), .Y(n_619) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_583), .B(n_598), .Y(n_643) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_583) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_638) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B(n_592), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_595), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g661 ( .A(n_595), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g700 ( .A(n_596), .B(n_618), .Y(n_700) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g743 ( .A(n_598), .B(n_653), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_599), .A2(n_716), .B1(n_718), .B2(n_721), .C(n_723), .Y(n_715) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g609 ( .A(n_601), .Y(n_609) );
OR2x2_ASAP7_75t_L g709 ( .A(n_601), .B(n_648), .Y(n_709) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_610), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_605), .A2(n_731), .B1(n_735), .B2(n_738), .Y(n_730) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
AND2x4_ASAP7_75t_L g654 ( .A(n_606), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g766 ( .A(n_606), .B(n_684), .Y(n_766) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g614 ( .A(n_608), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g630 ( .A(n_608), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g689 ( .A(n_608), .B(n_626), .Y(n_689) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_608), .Y(n_706) );
INVx1_ASAP7_75t_L g720 ( .A(n_608), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_608), .B(n_633), .Y(n_763) );
AND2x4_ASAP7_75t_L g670 ( .A(n_609), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g668 ( .A(n_611), .Y(n_668) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_612), .B(n_653), .Y(n_652) );
NAND2x1_ASAP7_75t_L g772 ( .A(n_612), .B(n_674), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B1(n_620), .B2(n_622), .Y(n_613) );
AND2x2_ASAP7_75t_L g639 ( .A(n_614), .B(n_632), .Y(n_639) );
INVx1_ASAP7_75t_L g680 ( .A(n_614), .Y(n_680) );
AND2x2_ASAP7_75t_L g787 ( .A(n_614), .B(n_648), .Y(n_787) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_618), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g760 ( .A(n_618), .Y(n_760) );
AND2x2_ASAP7_75t_L g777 ( .A(n_618), .B(n_637), .Y(n_777) );
AND2x2_ASAP7_75t_L g793 ( .A(n_618), .B(n_743), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_619), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g716 ( .A(n_619), .B(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_619), .A2(n_709), .B1(n_724), .B2(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g679 ( .A(n_621), .Y(n_679) );
AND2x2_ASAP7_75t_L g710 ( .A(n_621), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_621), .B(n_717), .Y(n_739) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g745 ( .A(n_625), .B(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_625), .A2(n_649), .B1(n_754), .B2(n_756), .Y(n_753) );
INVx3_ASAP7_75t_L g648 ( .A(n_626), .Y(n_648) );
AND2x2_ASAP7_75t_L g780 ( .A(n_626), .B(n_633), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_644), .Y(n_627) );
AOI32xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_634), .A3(n_637), .B1(n_639), .B2(n_640), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_631), .Y(n_726) );
INVx1_ASAP7_75t_L g751 ( .A(n_631), .Y(n_751) );
INVx3_ASAP7_75t_L g707 ( .A(n_632), .Y(n_707) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g782 ( .A1(n_635), .A2(n_783), .B1(n_784), .B2(n_785), .C(n_786), .Y(n_782) );
BUFx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g759 ( .A(n_637), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g795 ( .A(n_637), .B(n_756), .Y(n_795) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g653 ( .A(n_638), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_640), .B(n_668), .Y(n_667) );
AO22x1_ASAP7_75t_L g697 ( .A1(n_640), .A2(n_698), .B1(n_700), .B2(n_701), .Y(n_697) );
NAND2x1p5_ASAP7_75t_L g801 ( .A(n_640), .B(n_668), .Y(n_801) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g717 ( .A(n_641), .Y(n_717) );
INVx1_ASAP7_75t_L g727 ( .A(n_641), .Y(n_727) );
AND2x2_ASAP7_75t_L g647 ( .A(n_642), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_643), .Y(n_729) );
INVx1_ASAP7_75t_L g769 ( .A(n_643), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B(n_649), .C(n_654), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2x1p5_ASAP7_75t_L g756 ( .A(n_646), .B(n_676), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_647), .B(n_706), .Y(n_783) );
AOI31xp33_ASAP7_75t_L g666 ( .A1(n_648), .A2(n_667), .A3(n_669), .B(n_672), .Y(n_666) );
INVx4_ASAP7_75t_L g725 ( .A(n_648), .Y(n_725) );
OR2x2_ASAP7_75t_L g762 ( .A(n_648), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AND2x4_ASAP7_75t_L g664 ( .A(n_653), .B(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_655), .Y(n_660) );
AND2x2_ASAP7_75t_L g691 ( .A(n_655), .B(n_689), .Y(n_691) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_658), .B(n_666), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g784 ( .A(n_661), .Y(n_784) );
INVx1_ASAP7_75t_L g692 ( .A(n_662), .Y(n_692) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g722 ( .A(n_663), .Y(n_722) );
AND2x2_ASAP7_75t_L g721 ( .A(n_664), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .A3(n_681), .B1(n_685), .B2(n_688), .C1(n_690), .C2(n_692), .Y(n_678) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI211x1_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_697), .C(n_703), .Y(n_693) );
INVx1_ASAP7_75t_L g798 ( .A(n_694), .Y(n_798) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g752 ( .A(n_696), .Y(n_752) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OA21x2_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_708), .B(n_710), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx2_ASAP7_75t_L g773 ( .A(n_707), .Y(n_773) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp33_ASAP7_75t_L g768 ( .A(n_711), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_781), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_748), .C(n_764), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_730), .C(n_740), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_717), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI21xp33_ASAP7_75t_L g776 ( .A1(n_721), .A2(n_777), .B(n_778), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_725), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_725), .B(n_775), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_726), .B(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_727), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_737), .A2(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_744), .B(n_745), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_753), .C(n_757), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_SL g767 ( .A(n_759), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_763), .Y(n_785) );
OAI211xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B(n_770), .C(n_776), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_775), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g796 ( .A(n_775), .Y(n_796) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g792 ( .A(n_780), .Y(n_792) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_790), .C(n_797), .Y(n_781) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AOI21xp33_ASAP7_75t_SL g790 ( .A1(n_791), .A2(n_794), .B(n_796), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AOI21xp33_ASAP7_75t_R g797 ( .A1(n_798), .A2(n_799), .B(n_801), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx6_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx10_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OR2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_816), .Y(n_811) );
INVxp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
BUFx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
endmodule