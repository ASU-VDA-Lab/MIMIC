module real_aes_1949_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_0), .B(n_492), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_1), .A2(n_491), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_2), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_3), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_4), .B(n_209), .Y(n_562) );
INVx1_ASAP7_75t_L g137 ( .A(n_5), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_6), .B(n_146), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_7), .B(n_209), .Y(n_529) );
INVx1_ASAP7_75t_L g243 ( .A(n_8), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_9), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_10), .Y(n_257) );
NAND2xp33_ASAP7_75t_L g539 ( .A(n_11), .B(n_206), .Y(n_539) );
INVx2_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
AOI221x1_ASAP7_75t_L g490 ( .A1(n_13), .A2(n_25), .B1(n_491), .B2(n_492), .C(n_493), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
AND3x1_ASAP7_75t_L g788 ( .A(n_14), .B(n_40), .C(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_15), .B(n_492), .Y(n_535) );
INVx1_ASAP7_75t_L g207 ( .A(n_16), .Y(n_207) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_17), .A2(n_168), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_18), .B(n_184), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_19), .B(n_209), .Y(n_546) );
AO21x1_ASAP7_75t_L g557 ( .A1(n_20), .A2(n_492), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_L g204 ( .A(n_22), .Y(n_204) );
INVx1_ASAP7_75t_SL g190 ( .A(n_23), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_24), .B(n_157), .Y(n_156) );
AOI33xp33_ASAP7_75t_L g223 ( .A1(n_26), .A2(n_54), .A3(n_134), .B1(n_152), .B2(n_224), .B3(n_225), .Y(n_223) );
NAND2x1_ASAP7_75t_L g502 ( .A(n_27), .B(n_209), .Y(n_502) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_28), .B(n_206), .Y(n_528) );
INVx1_ASAP7_75t_L g251 ( .A(n_29), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_30), .Y(n_104) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_31), .A2(n_85), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g147 ( .A(n_31), .B(n_85), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_32), .B(n_178), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_33), .B(n_206), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g116 ( .A1(n_34), .A2(n_117), .B1(n_762), .B2(n_763), .C(n_768), .Y(n_116) );
INVx1_ASAP7_75t_L g762 ( .A(n_34), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_35), .B(n_209), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_36), .A2(n_766), .B1(n_781), .B2(n_782), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_36), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_37), .B(n_206), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_38), .A2(n_491), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g140 ( .A(n_39), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g151 ( .A(n_39), .Y(n_151) );
AND2x2_ASAP7_75t_L g166 ( .A(n_39), .B(n_137), .Y(n_166) );
OR2x6_ASAP7_75t_L g112 ( .A(n_40), .B(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_41), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_42), .B(n_492), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_43), .B(n_178), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_44), .A2(n_131), .B1(n_143), .B2(n_146), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_45), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_46), .B(n_157), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_47), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_48), .B(n_206), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_49), .B(n_168), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_50), .B(n_157), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_51), .A2(n_491), .B(n_527), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_52), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_53), .B(n_206), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_55), .B(n_157), .Y(n_235) );
INVx1_ASAP7_75t_L g135 ( .A(n_56), .Y(n_135) );
INVx1_ASAP7_75t_L g159 ( .A(n_56), .Y(n_159) );
AND2x2_ASAP7_75t_L g236 ( .A(n_57), .B(n_184), .Y(n_236) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_58), .A2(n_74), .B1(n_149), .B2(n_178), .C(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_59), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_60), .B(n_209), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_61), .B(n_143), .Y(n_259) );
AOI21xp5_ASAP7_75t_SL g173 ( .A1(n_62), .A2(n_149), .B(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_63), .A2(n_491), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g200 ( .A(n_64), .Y(n_200) );
AO21x1_ASAP7_75t_L g559 ( .A1(n_65), .A2(n_491), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_66), .B(n_492), .Y(n_519) );
INVx1_ASAP7_75t_L g234 ( .A(n_67), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_68), .B(n_492), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_69), .A2(n_149), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g513 ( .A(n_70), .B(n_185), .Y(n_513) );
INVx1_ASAP7_75t_L g141 ( .A(n_71), .Y(n_141) );
INVx1_ASAP7_75t_L g161 ( .A(n_71), .Y(n_161) );
AND2x2_ASAP7_75t_L g531 ( .A(n_72), .B(n_171), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_73), .B(n_178), .Y(n_226) );
AND2x2_ASAP7_75t_L g192 ( .A(n_75), .B(n_171), .Y(n_192) );
INVx1_ASAP7_75t_L g201 ( .A(n_76), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_77), .A2(n_149), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_78), .A2(n_149), .B(n_155), .C(n_167), .Y(n_148) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
AND2x2_ASAP7_75t_L g517 ( .A(n_80), .B(n_171), .Y(n_517) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_81), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_82), .B(n_492), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_83), .A2(n_149), .B1(n_221), .B2(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g558 ( .A(n_84), .B(n_146), .Y(n_558) );
AND2x2_ASAP7_75t_L g505 ( .A(n_86), .B(n_171), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_87), .B(n_206), .Y(n_547) );
INVx1_ASAP7_75t_L g175 ( .A(n_88), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_89), .B(n_209), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_90), .B(n_206), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_91), .A2(n_491), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g227 ( .A(n_92), .B(n_171), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_93), .B(n_209), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_94), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_95), .Y(n_769) );
BUFx2_ASAP7_75t_L g775 ( .A(n_96), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_97), .A2(n_491), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_98), .B(n_157), .Y(n_176) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_784), .B(n_792), .Y(n_99) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_771), .B(n_776), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_116), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_103), .A2(n_780), .B(n_783), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g783 ( .A(n_107), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_SL g120 ( .A(n_110), .B(n_111), .Y(n_120) );
AND2x6_ASAP7_75t_SL g480 ( .A(n_110), .B(n_112), .Y(n_480) );
OR2x2_ASAP7_75t_L g770 ( .A(n_110), .B(n_112), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g787 ( .A(n_113), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_121), .B1(n_477), .B2(n_481), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
CKINVDCx11_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_120), .A2(n_764), .B1(n_766), .B2(n_767), .Y(n_763) );
INVxp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g765 ( .A(n_122), .Y(n_765) );
NAND4xp75_ASAP7_75t_L g122 ( .A(n_123), .B(n_328), .C(n_394), .D(n_457), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_291), .Y(n_123) );
OR3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_261), .C(n_288), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_193), .B(n_216), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_179), .Y(n_127) );
AND2x2_ASAP7_75t_L g391 ( .A(n_128), .B(n_361), .Y(n_391) );
INVx1_ASAP7_75t_L g464 ( .A(n_128), .Y(n_464) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_169), .Y(n_128) );
INVx2_ASAP7_75t_L g215 ( .A(n_129), .Y(n_215) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_129), .Y(n_279) );
AND2x2_ASAP7_75t_L g283 ( .A(n_129), .B(n_196), .Y(n_283) );
AND2x4_ASAP7_75t_L g299 ( .A(n_129), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g303 ( .A(n_129), .Y(n_303) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_148), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_138), .C(n_142), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g178 ( .A(n_133), .B(n_139), .Y(n_178) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
OR2x6_ASAP7_75t_L g164 ( .A(n_134), .B(n_153), .Y(n_164) );
INVxp33_ASAP7_75t_L g224 ( .A(n_134), .Y(n_224) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g154 ( .A(n_135), .B(n_137), .Y(n_154) );
AND2x4_ASAP7_75t_L g209 ( .A(n_135), .B(n_160), .Y(n_209) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g491 ( .A(n_140), .B(n_154), .Y(n_491) );
INVx2_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
AND2x6_ASAP7_75t_L g206 ( .A(n_141), .B(n_158), .Y(n_206) );
INVx4_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_143), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AND2x4_ASAP7_75t_L g146 ( .A(n_145), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_145), .B(n_147), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_146), .A2(n_173), .B(n_177), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_146), .B(n_165), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_146), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_SL g542 ( .A(n_146), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_146), .B(n_564), .Y(n_563) );
INVxp67_ASAP7_75t_L g258 ( .A(n_149), .Y(n_258) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NOR2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_162), .B(n_165), .Y(n_155) );
INVx1_ASAP7_75t_L g202 ( .A(n_157), .Y(n_202) );
AND2x4_ASAP7_75t_L g492 ( .A(n_157), .B(n_166), .Y(n_492) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_164), .A2(n_165), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_164), .A2(n_165), .B(n_190), .C(n_191), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_164), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_164), .A2(n_165), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_164), .A2(n_165), .B(n_243), .C(n_244), .Y(n_242) );
INVxp67_ASAP7_75t_L g249 ( .A(n_164), .Y(n_249) );
INVx1_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_165), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_165), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_165), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_165), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_165), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_165), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_165), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_165), .A2(n_561), .B(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_166), .Y(n_252) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_167), .A2(n_219), .B(n_227), .Y(n_218) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_167), .A2(n_219), .B(n_227), .Y(n_267) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_168), .A2(n_241), .B(n_245), .Y(n_240) );
AND2x2_ASAP7_75t_L g194 ( .A(n_169), .B(n_195), .Y(n_194) );
INVx4_ASAP7_75t_L g280 ( .A(n_169), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_169), .B(n_270), .Y(n_284) );
INVx2_ASAP7_75t_L g298 ( .A(n_169), .Y(n_298) );
AND2x4_ASAP7_75t_L g302 ( .A(n_169), .B(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_169), .Y(n_337) );
OR2x2_ASAP7_75t_L g343 ( .A(n_169), .B(n_182), .Y(n_343) );
NOR2x1_ASAP7_75t_SL g372 ( .A(n_169), .B(n_196), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_169), .B(n_446), .Y(n_474) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_172), .Y(n_169) );
INVx3_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_171), .A2(n_229), .B1(n_248), .B2(n_253), .Y(n_247) );
INVx1_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
AND2x2_ASAP7_75t_L g371 ( .A(n_179), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2x1_ASAP7_75t_L g405 ( .A(n_180), .B(n_195), .Y(n_405) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g212 ( .A(n_182), .Y(n_212) );
INVx2_ASAP7_75t_L g271 ( .A(n_182), .Y(n_271) );
AND2x2_ASAP7_75t_L g294 ( .A(n_182), .B(n_196), .Y(n_294) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_182), .Y(n_321) );
INVx1_ASAP7_75t_L g362 ( .A(n_182), .Y(n_362) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_192), .Y(n_182) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_183), .A2(n_525), .B(n_531), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_184), .A2(n_490), .B(n_496), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_184), .A2(n_519), .B(n_520), .Y(n_518) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_184), .A2(n_490), .B(n_496), .Y(n_598) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_211), .Y(n_193) );
AND2x2_ASAP7_75t_L g374 ( .A(n_194), .B(n_269), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_195), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g441 ( .A(n_195), .Y(n_441) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g300 ( .A(n_196), .Y(n_300) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_203), .B(n_210), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_202), .B(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B1(n_207), .B2(n_208), .Y(n_203) );
INVxp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_211), .A2(n_378), .B(n_382), .C(n_388), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_213), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_SL g424 ( .A(n_213), .Y(n_424) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g346 ( .A(n_215), .B(n_300), .Y(n_346) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_237), .Y(n_216) );
AOI32xp33_ASAP7_75t_L g382 ( .A1(n_217), .A2(n_366), .A3(n_383), .B1(n_384), .B2(n_386), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
INVx2_ASAP7_75t_L g308 ( .A(n_218), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_218), .B(n_240), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_220), .B(n_226), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_228), .B(n_246), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_228), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_228), .Y(n_438) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_236), .Y(n_228) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_229), .A2(n_230), .B(n_236), .Y(n_266) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_229), .A2(n_499), .B(n_505), .Y(n_498) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_229), .A2(n_507), .B(n_513), .Y(n_506) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_229), .A2(n_507), .B(n_513), .Y(n_565) );
AO21x2_ASAP7_75t_L g590 ( .A1(n_229), .A2(n_499), .B(n_505), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
OR2x2_ASAP7_75t_L g339 ( .A(n_237), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g290 ( .A(n_238), .B(n_264), .Y(n_290) );
AND2x2_ASAP7_75t_L g439 ( .A(n_238), .B(n_437), .Y(n_439) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_246), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g276 ( .A(n_240), .Y(n_276) );
AND2x4_ASAP7_75t_L g315 ( .A(n_240), .B(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_L g349 ( .A(n_240), .Y(n_349) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_240), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_240), .B(n_246), .Y(n_366) );
INVx1_ASAP7_75t_L g450 ( .A(n_240), .Y(n_450) );
INVx2_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
INVx1_ASAP7_75t_L g314 ( .A(n_246), .Y(n_314) );
INVx1_ASAP7_75t_L g381 ( .A(n_246), .Y(n_381) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_258), .B1(n_259), .B2(n_260), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI32xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_272), .A3(n_277), .B1(n_281), .B2(n_285), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_263), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_264), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_264), .B(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g390 ( .A(n_264), .Y(n_390) );
AND2x2_ASAP7_75t_L g471 ( .A(n_264), .B(n_313), .Y(n_471) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g385 ( .A(n_266), .B(n_308), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_266), .B(n_287), .Y(n_407) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_266), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
INVx1_ASAP7_75t_L g340 ( .A(n_267), .Y(n_340) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_287), .Y(n_355) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g383 ( .A(n_269), .B(n_372), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_269), .B(n_302), .Y(n_453) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_270), .Y(n_422) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_271), .Y(n_404) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g305 ( .A(n_274), .B(n_306), .Y(n_305) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_274), .B(n_390), .Y(n_389) );
NOR2xp67_ASAP7_75t_SL g476 ( .A(n_274), .B(n_414), .Y(n_476) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g333 ( .A(n_276), .B(n_287), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_277), .B(n_343), .Y(n_401) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_278), .B(n_294), .Y(n_367) );
AND2x4_ASAP7_75t_SL g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_280), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g432 ( .A(n_280), .B(n_303), .Y(n_432) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_280), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_281), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
OR2x2_ASAP7_75t_L g403 ( .A(n_282), .B(n_404), .Y(n_403) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_282), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g392 ( .A(n_283), .B(n_337), .Y(n_392) );
INVxp33_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_286), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g466 ( .A(n_286), .B(n_348), .Y(n_466) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_309), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_295), .B(n_304), .Y(n_292) );
AND2x2_ASAP7_75t_L g427 ( .A(n_294), .B(n_302), .Y(n_427) );
NAND2xp33_ASAP7_75t_R g295 ( .A(n_296), .B(n_301), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g469 ( .A(n_298), .Y(n_469) );
INVx4_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
INVx1_ASAP7_75t_L g446 ( .A(n_300), .Y(n_446) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g440 ( .A(n_302), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_302), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_305), .A2(n_370), .B1(n_474), .B2(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g334 ( .A(n_308), .B(n_320), .Y(n_334) );
AND2x2_ASAP7_75t_L g348 ( .A(n_308), .B(n_349), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_317), .B(n_322), .C(n_325), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g396 ( .A(n_312), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_313), .Y(n_324) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g384 ( .A(n_314), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g393 ( .A(n_314), .B(n_315), .Y(n_393) );
INVx1_ASAP7_75t_L g425 ( .A(n_314), .Y(n_425) );
AND2x4_ASAP7_75t_L g406 ( .A(n_315), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_315), .B(n_319), .Y(n_428) );
AND2x2_ASAP7_75t_L g436 ( .A(n_315), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g411 ( .A(n_319), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_319), .B(n_333), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_319), .B(n_366), .Y(n_416) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_320), .B(n_381), .Y(n_430) );
AND2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_346), .Y(n_358) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g454 ( .A(n_324), .B(n_334), .Y(n_454) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_326), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g338 ( .A(n_327), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_327), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_368), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_352), .Y(n_329) );
OAI222xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_339), .B2(n_341), .C1(n_344), .C2(n_347), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_337), .B(n_346), .Y(n_345) );
OR2x6_ASAP7_75t_L g417 ( .A(n_337), .B(n_387), .Y(n_417) );
NAND5xp2_ASAP7_75t_L g420 ( .A(n_337), .B(n_340), .C(n_356), .D(n_421), .E(n_423), .Y(n_420) );
NAND2x1_ASAP7_75t_L g456 ( .A(n_338), .B(n_342), .Y(n_456) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_343), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_345), .A2(n_436), .B1(n_439), .B2(n_440), .Y(n_435) );
INVx2_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_346), .B(n_362), .Y(n_399) );
INVx3_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g379 ( .A(n_348), .B(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g412 ( .A(n_348), .Y(n_412) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g375 ( .A(n_351), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_364), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B(n_359), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g363 ( .A(n_355), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_358), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_SL g445 ( .A(n_362), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_377), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_388) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_418), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .C(n_408), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OA21x2_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B(n_406), .Y(n_400) );
NAND2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_415), .B(n_417), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_412), .A2(n_452), .B1(n_454), .B2(n_455), .Y(n_451) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_442), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .C(n_433), .D(n_435), .Y(n_419) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g431 ( .A(n_422), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_429), .B2(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_431), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_447), .B(n_451), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_470), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx4_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
CKINVDCx11_ASAP7_75t_R g767 ( .A(n_480), .Y(n_767) );
INVx3_ASAP7_75t_L g766 ( .A(n_481), .Y(n_766) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_674), .Y(n_481) );
AND4x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_586), .C(n_613), .D(n_648), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_514), .B1(n_551), .B2(n_566), .C(n_570), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_486), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g627 ( .A(n_487), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_637), .Y(n_682) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g585 ( .A(n_488), .B(n_506), .Y(n_585) );
AND2x4_ASAP7_75t_L g621 ( .A(n_488), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g635 ( .A(n_488), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g552 ( .A(n_489), .Y(n_552) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_489), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_SL g579 ( .A1(n_497), .A2(n_552), .B(n_580), .C(n_584), .Y(n_579) );
AND2x2_ASAP7_75t_L g600 ( .A(n_497), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_497), .B(n_552), .Y(n_740) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_506), .Y(n_497) );
INVx2_ASAP7_75t_L g620 ( .A(n_498), .Y(n_620) );
BUFx3_ASAP7_75t_L g636 ( .A(n_498), .Y(n_636) );
INVxp67_ASAP7_75t_L g640 ( .A(n_498), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .Y(n_499) );
INVx2_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_506), .B(n_598), .Y(n_625) );
AND2x2_ASAP7_75t_L g651 ( .A(n_506), .B(n_620), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_514), .A2(n_649), .B(n_652), .C(n_662), .Y(n_648) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_532), .Y(n_514) );
OAI321xp33_ASAP7_75t_L g623 ( .A1(n_515), .A2(n_571), .A3(n_624), .B1(n_626), .B2(n_627), .C(n_629), .Y(n_623) );
AND2x2_ASAP7_75t_L g744 ( .A(n_515), .B(n_719), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_515), .Y(n_747) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
INVx5_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_516), .B(n_583), .Y(n_582) );
NOR2x1_ASAP7_75t_SL g614 ( .A(n_516), .B(n_615), .Y(n_614) );
BUFx2_ASAP7_75t_L g659 ( .A(n_516), .Y(n_659) );
AND2x2_ASAP7_75t_L g761 ( .A(n_516), .B(n_533), .Y(n_761) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g568 ( .A(n_524), .B(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
INVx4_ASAP7_75t_L g583 ( .A(n_524), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g626 ( .A(n_532), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_R g729 ( .A1(n_532), .A2(n_568), .B(n_600), .C(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g749 ( .A(n_532), .B(n_574), .Y(n_749) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_540), .Y(n_532) );
INVx1_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
INVx2_ASAP7_75t_L g573 ( .A(n_533), .Y(n_573) );
OR2x2_ASAP7_75t_L g592 ( .A(n_533), .B(n_583), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_533), .B(n_615), .Y(n_661) );
BUFx3_ASAP7_75t_L g668 ( .A(n_533), .Y(n_668) );
INVx1_ASAP7_75t_L g631 ( .A(n_540), .Y(n_631) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_540), .Y(n_644) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g577 ( .A(n_541), .Y(n_577) );
INVx1_ASAP7_75t_L g686 ( .A(n_541), .Y(n_686) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_542), .B(n_550), .Y(n_549) );
AO21x2_ASAP7_75t_L g615 ( .A1(n_542), .A2(n_543), .B(n_549), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
AND2x2_ASAP7_75t_L g587 ( .A(n_551), .B(n_588), .Y(n_587) );
OAI31xp33_ASAP7_75t_L g738 ( .A1(n_551), .A2(n_739), .A3(n_741), .B(n_744), .Y(n_738) );
INVx1_ASAP7_75t_SL g756 ( .A(n_551), .Y(n_756) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g570 ( .A1(n_552), .A2(n_571), .B(n_579), .Y(n_570) );
NAND2x1_ASAP7_75t_L g650 ( .A(n_552), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g679 ( .A(n_552), .Y(n_679) );
INVx2_ASAP7_75t_L g628 ( .A(n_553), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_553), .B(n_611), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_553), .B(n_610), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g728 ( .A(n_553), .B(n_679), .Y(n_728) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_565), .Y(n_553) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_554), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g608 ( .A(n_554), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g637 ( .A(n_554), .B(n_619), .Y(n_637) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g622 ( .A(n_556), .Y(n_622) );
OAI21x1_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_559), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g564 ( .A(n_558), .Y(n_564) );
INVx2_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_565), .Y(n_669) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g605 ( .A(n_567), .Y(n_605) );
AND2x2_ASAP7_75t_L g684 ( .A(n_567), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_589), .Y(n_595) );
INVx2_ASAP7_75t_SL g643 ( .A(n_568), .Y(n_643) );
INVx4_ASAP7_75t_L g574 ( .A(n_569), .Y(n_574) );
AND2x2_ASAP7_75t_L g672 ( .A(n_569), .B(n_615), .Y(n_672) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_569), .B(n_685), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g707 ( .A(n_569), .B(n_583), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_571), .Y(n_713) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
OR2x2_ASAP7_75t_L g645 ( .A(n_572), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
OR2x2_ASAP7_75t_L g697 ( .A(n_573), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g727 ( .A(n_573), .B(n_615), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_574), .B(n_577), .Y(n_603) );
AND2x2_ASAP7_75t_L g695 ( .A(n_574), .B(n_685), .Y(n_695) );
AND2x4_ASAP7_75t_L g757 ( .A(n_574), .B(n_636), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx2_ASAP7_75t_L g581 ( .A(n_576), .Y(n_581) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp67_ASAP7_75t_SL g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OAI322xp33_ASAP7_75t_SL g593 ( .A1(n_581), .A2(n_594), .A3(n_596), .B1(n_599), .B2(n_602), .C1(n_604), .C2(n_606), .Y(n_593) );
INVx1_ASAP7_75t_L g751 ( .A(n_581), .Y(n_751) );
OR2x2_ASAP7_75t_L g604 ( .A(n_582), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g630 ( .A(n_583), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_583), .B(n_631), .Y(n_646) );
INVx2_ASAP7_75t_L g673 ( .A(n_583), .Y(n_673) );
AND2x4_ASAP7_75t_L g685 ( .A(n_583), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_585), .B(n_601), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_591), .B(n_593), .Y(n_586) );
AND2x2_ASAP7_75t_L g654 ( .A(n_588), .B(n_621), .Y(n_654) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_589), .B(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g612 ( .A(n_590), .Y(n_612) );
AND2x4_ASAP7_75t_SL g694 ( .A(n_590), .B(n_609), .Y(n_694) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g602 ( .A(n_592), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_595), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g730 ( .A(n_597), .B(n_694), .Y(n_730) );
NOR4xp25_ASAP7_75t_L g734 ( .A(n_597), .B(n_611), .C(n_651), .D(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g611 ( .A(n_598), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g647 ( .A(n_598), .B(n_622), .Y(n_647) );
AND2x4_ASAP7_75t_L g711 ( .A(n_598), .B(n_622), .Y(n_711) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_601), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
OR2x2_ASAP7_75t_L g700 ( .A(n_608), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g754 ( .A(n_608), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_609), .B(n_621), .Y(n_655) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AOI211xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_616), .B(n_623), .C(n_638), .Y(n_613) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_619), .B(n_622), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_620), .B(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g702 ( .A(n_620), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_621), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g717 ( .A(n_621), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_633), .Y(n_629) );
AND2x4_ASAP7_75t_L g666 ( .A(n_630), .B(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g760 ( .A(n_630), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_SL g664 ( .A(n_636), .Y(n_664) );
AND2x2_ASAP7_75t_L g723 ( .A(n_637), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
O2A1O1Ixp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_641), .B(n_645), .C(n_647), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_639), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g715 ( .A(n_640), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g736 ( .A(n_640), .B(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OR2x2_ASAP7_75t_L g725 ( .A(n_643), .B(n_667), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_646), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_652) );
INVx1_ASAP7_75t_SL g743 ( .A(n_647), .Y(n_743) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_658), .B(n_667), .Y(n_709) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_661), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B1(n_669), .B2(n_670), .Y(n_662) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI21xp5_ASAP7_75t_SL g676 ( .A1(n_667), .A2(n_677), .B(n_680), .Y(n_676) );
AND2x2_ASAP7_75t_L g705 ( .A(n_667), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND3x2_ASAP7_75t_L g671 ( .A(n_668), .B(n_672), .C(n_673), .Y(n_671) );
AND2x2_ASAP7_75t_L g733 ( .A(n_668), .B(n_690), .Y(n_733) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g718 ( .A(n_673), .B(n_719), .Y(n_718) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_675), .B(n_731), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_691), .C(n_712), .D(n_729), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_687), .B2(n_689), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_683), .A2(n_697), .B1(n_717), .B2(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g698 ( .A(n_685), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_687), .A2(n_710), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx3_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B1(n_696), .B2(n_699), .C(n_703), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_706), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_706), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_718), .B2(n_720), .C(n_721), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_717), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B1(n_726), .B2(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g746 ( .A1(n_727), .A2(n_747), .B(n_748), .C(n_750), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B(n_738), .C(n_745), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_752), .B1(n_755), .B2(n_757), .C(n_758), .Y(n_745) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g782 ( .A(n_766), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
BUFx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_775), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_786), .Y(n_795) );
AND2x2_ASAP7_75t_SL g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
endmodule