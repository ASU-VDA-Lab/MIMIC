module fake_jpeg_8526_n_267 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_14),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_58),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_30),
.B1(n_20),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_62),
.B1(n_20),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_20),
.B2(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_41),
.Y(n_81)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_86),
.Y(n_111)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_41),
.C(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_90),
.B(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_31),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_31),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_27),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g88 ( 
.A(n_58),
.Y(n_88)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_27),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_34),
.C(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_84),
.Y(n_127)
);

CKINVDCx11_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_64),
.B1(n_61),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_116),
.CON(n_130),
.SN(n_130)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_61),
.B1(n_64),
.B2(n_22),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_61),
.B1(n_66),
.B2(n_22),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_108),
.B1(n_86),
.B2(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_79),
.B(n_90),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_71),
.B(n_79),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_125),
.B(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_124),
.Y(n_163)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_75),
.C(n_70),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_136),
.C(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_131),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_69),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_89),
.C(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_56),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_95),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_128),
.B1(n_118),
.B2(n_107),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_45),
.B1(n_76),
.B2(n_2),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_119),
.B(n_138),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_149),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_107),
.B1(n_101),
.B2(n_120),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_166),
.B1(n_109),
.B2(n_103),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_164),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_111),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_141),
.C(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_107),
.B1(n_100),
.B2(n_95),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_109),
.B1(n_45),
.B2(n_73),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_102),
.B(n_108),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_106),
.B(n_104),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_162),
.B(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_167),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_25),
.B(n_22),
.Y(n_165)
);

AO22x2_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_115),
.B1(n_29),
.B2(n_34),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_169),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_125),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_173),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_137),
.B1(n_122),
.B2(n_31),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_182),
.C(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_181),
.B1(n_184),
.B2(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_46),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_109),
.B1(n_76),
.B2(n_73),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_46),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_147),
.C(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_143),
.B1(n_162),
.B2(n_153),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_76),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_165),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_159),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_197),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_171),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_145),
.B1(n_144),
.B2(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_175),
.C(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_207),
.C(n_209),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_210),
.B1(n_188),
.B2(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_176),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_149),
.C(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_197),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_174),
.C(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.C(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_181),
.C(n_190),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_221),
.Y(n_229)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_173),
.C(n_187),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_201),
.B1(n_208),
.B2(n_210),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_186),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_185),
.C(n_4),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_234),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_232),
.B1(n_223),
.B2(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_202),
.B1(n_192),
.B2(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_196),
.B1(n_185),
.B2(n_156),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_235),
.B1(n_3),
.B2(n_4),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_185),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_216),
.B1(n_213),
.B2(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_5),
.C(n_6),
.Y(n_246)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_242),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_214),
.B(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_3),
.C(n_5),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_230),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_227),
.B(n_232),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_252),
.B(n_246),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_237),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_238),
.C(n_7),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_235),
.B(n_7),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_8),
.A3(n_10),
.B1(n_13),
.B2(n_15),
.C1(n_16),
.C2(n_248),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_255),
.A2(n_253),
.B1(n_9),
.B2(n_10),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_8),
.C(n_13),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_13),
.B(n_16),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_264),
.B(n_262),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_261),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_259),
.Y(n_267)
);


endmodule