module real_jpeg_4455_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_1),
.A2(n_33),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_33),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_93),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_1),
.A2(n_237),
.B(n_309),
.C(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_1),
.B(n_333),
.C(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_1),
.B(n_117),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_1),
.B(n_157),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_1),
.B(n_61),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_83),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_2),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_179),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_2),
.A2(n_179),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_2),
.A2(n_179),
.B1(n_343),
.B2(n_345),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_5),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_68),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_6),
.A2(n_68),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_6),
.A2(n_68),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_44),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_44),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_11),
.Y(n_333)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_208),
.B1(n_401),
.B2(n_402),
.Y(n_13)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_14),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_206),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_184),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_16),
.B(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_109),
.C(n_151),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_17),
.A2(n_109),
.B1(n_110),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_74),
.B2(n_75),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_18),
.A2(n_76),
.B(n_78),
.Y(n_205)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_20),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_20),
.A2(n_37),
.B1(n_76),
.B2(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_20),
.B(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_20),
.A2(n_76),
.B1(n_308),
.B2(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_29),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_21),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_21),
.B(n_29),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_21),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_21),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_24),
.Y(n_165)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_33),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_33),
.B(n_107),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_33),
.A2(n_311),
.B(n_314),
.Y(n_310)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_37),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_47),
.B(n_66),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_38),
.A2(n_147),
.B(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_43),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_47),
.A2(n_141),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_48),
.B(n_67),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_48),
.B(n_142),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_48),
.B(n_321),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_61),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_59),
.A2(n_119),
.B1(n_122),
.B2(n_124),
.Y(n_118)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_59),
.Y(n_323)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_61),
.B(n_321),
.Y(n_337)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g259 ( 
.A(n_66),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_66),
.B(n_320),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_70),
.B(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_73),
.Y(n_316)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_101),
.B(n_102),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_80),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_80),
.B(n_103),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_80),
.B(n_191),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_93),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_91),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_86),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_93),
.B(n_103),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_93),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_93),
.B(n_178),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_94),
.Y(n_233)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_97),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_99),
.Y(n_232)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_106),
.Y(n_234)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_139),
.B(n_150),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_139),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B(n_126),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_112),
.A2(n_170),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_117),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_117),
.A2(n_170),
.B(n_171),
.Y(n_277)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_118),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_120),
.Y(n_313)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_121),
.Y(n_309)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_148),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_140),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_149),
.B(n_337),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_186),
.B1(n_187),
.B2(n_204),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_151),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_167),
.C(n_175),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_152),
.A2(n_153),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_166),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_154),
.B(n_166),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_155),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_156),
.A2(n_160),
.B(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_159),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_161),
.B(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_162),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_164),
.Y(n_344)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_167),
.B(n_175),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_169),
.B(n_219),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_170),
.B(n_220),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_171),
.Y(n_268)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_190),
.Y(n_264)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_231),
.A3(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_205),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_197),
.B2(n_198),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_200),
.B1(n_217),
.B2(n_227),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_214),
.C(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_393),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_283),
.C(n_298),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_269),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_253),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_212),
.B(n_253),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_228),
.C(n_244),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_213),
.B(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_215),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_228),
.A2(n_229),
.B1(n_244),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_239),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_239),
.Y(n_262)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

INVx6_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_251),
.B(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_245),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_249),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_250),
.B(n_357),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_251),
.B(n_341),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_264),
.C(n_265),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_269),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_282),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_270),
.B(n_282),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_295),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_284),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_285),
.B(n_292),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_289),
.CI(n_291),
.CON(n_296),
.SN(n_296)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_295),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_296),
.B(n_297),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_296),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_325),
.B(n_392),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_300),
.B(n_303),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.C(n_317),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_307),
.A2(n_317),
.B1(n_318),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_386),
.B(n_391),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_376),
.B(n_385),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_351),
.B(n_375),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_338),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_338),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_336),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_330),
.A2(n_331),
.B1(n_336),
.B2(n_354),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_349),
.C(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_362),
.B(n_374),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_355),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_370),
.B(n_373),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_372),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_379),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.C(n_383),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_390),
.Y(n_391)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_395),
.B(n_398),
.C(n_399),
.D(n_400),
.Y(n_393)
);


endmodule