module fake_jpeg_5025_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_10),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_25),
.C(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_11),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_22),
.B1(n_20),
.B2(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_11),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.C(n_11),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_19),
.C(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_30),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.C(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

NAND2xp67_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_16),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_16),
.C(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.C(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_27),
.C(n_12),
.Y(n_66)
);

OAI322xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_50),
.A3(n_56),
.B1(n_55),
.B2(n_53),
.C1(n_19),
.C2(n_12),
.Y(n_63)
);

AOI31xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_57),
.A3(n_12),
.B(n_13),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_66),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_57),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_69),
.Y(n_72)
);

AOI31xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_13),
.A3(n_2),
.B(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_13),
.B1(n_8),
.B2(n_3),
.Y(n_69)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_13),
.C(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_72),
.B1(n_73),
.B2(n_6),
.Y(n_76)
);

AOI211xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_75),
.B(n_4),
.C(n_7),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_1),
.Y(n_78)
);


endmodule