module fake_jpeg_6132_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_21),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_57),
.B1(n_26),
.B2(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_17),
.B1(n_29),
.B2(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_30),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_17),
.B1(n_33),
.B2(n_29),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_72),
.B(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_62),
.B1(n_43),
.B2(n_27),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_33),
.B1(n_39),
.B2(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_44),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_37),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_20),
.Y(n_90)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_35),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_28),
.B(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_59),
.B(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_28),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_57),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_63),
.B(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_95),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_87),
.B1(n_89),
.B2(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_18),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_109),
.B1(n_37),
.B2(n_24),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_30),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_76),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_86),
.C(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_114),
.B1(n_85),
.B2(n_81),
.Y(n_117)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_109)
);

AOI22x1_ASAP7_75t_R g124 ( 
.A1(n_112),
.A2(n_58),
.B1(n_37),
.B2(n_95),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_52),
.B1(n_67),
.B2(n_63),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.C(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_119),
.C(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_88),
.B1(n_83),
.B2(n_79),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_117),
.B1(n_127),
.B2(n_120),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_90),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_20),
.C(n_22),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_129),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_17),
.B1(n_54),
.B2(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_103),
.Y(n_136)
);

FAx1_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_30),
.CI(n_24),
.CON(n_129),
.SN(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_98),
.A3(n_107),
.B1(n_97),
.B2(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_136),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_146),
.B(n_20),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_144),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_97),
.A3(n_105),
.B1(n_113),
.B2(n_102),
.C(n_24),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_25),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_105),
.B1(n_104),
.B2(n_24),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_121),
.C(n_22),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_119),
.B1(n_115),
.B2(n_130),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_141),
.B(n_135),
.C(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_160),
.C(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_80),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_146),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_22),
.B(n_25),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_80),
.C(n_20),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_22),
.C(n_23),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_22),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_170),
.B(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_13),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.C(n_22),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_134),
.C(n_147),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_146),
.B1(n_142),
.B2(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_14),
.B1(n_13),
.B2(n_15),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_25),
.B1(n_23),
.B2(n_15),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_161),
.B1(n_159),
.B2(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_160),
.B(n_14),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_180),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_25),
.C(n_23),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_1),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_3),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_5),
.C(n_7),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_3),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_188),
.B(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_173),
.B1(n_174),
.B2(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_191),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_177),
.C(n_5),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_8),
.B(n_10),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_4),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_194),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_8),
.B(n_9),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_8),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_200),
.B(n_11),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_190),
.A3(n_186),
.B1(n_15),
.B2(n_23),
.C1(n_12),
.C2(n_11),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_196),
.B1(n_12),
.B2(n_11),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);


endmodule