module fake_netlist_1_5789_n_500 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_500);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_500;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_393;
wire n_135;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_69;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g63 ( .A(n_1), .Y(n_63) );
INVx2_ASAP7_75t_L g64 ( .A(n_27), .Y(n_64) );
INVxp33_ASAP7_75t_L g65 ( .A(n_39), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_49), .Y(n_66) );
CKINVDCx16_ASAP7_75t_R g67 ( .A(n_41), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_48), .Y(n_68) );
INVxp67_ASAP7_75t_L g69 ( .A(n_36), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_28), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_53), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_7), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_22), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_55), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_38), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_61), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_54), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_44), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_52), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_15), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_37), .B(n_18), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_42), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_6), .B(n_16), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_47), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_29), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_25), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_60), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_0), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_11), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_51), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_6), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_66), .Y(n_98) );
INVx2_ASAP7_75t_SL g99 ( .A(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_96), .B(n_0), .Y(n_101) );
AND2x4_ASAP7_75t_L g102 ( .A(n_87), .B(n_1), .Y(n_102) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_68), .B(n_35), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_81), .B(n_65), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_67), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_67), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_83), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_68), .A2(n_2), .B(n_3), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_63), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_63), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_94), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_70), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_88), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_91), .Y(n_118) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_64), .A2(n_34), .B(n_59), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_71), .Y(n_121) );
INVx4_ASAP7_75t_L g122 ( .A(n_102), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_113), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_113), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_113), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_113), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_99), .B(n_92), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_119), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g130 ( .A(n_103), .B(n_85), .Y(n_130) );
INVx2_ASAP7_75t_SL g131 ( .A(n_105), .Y(n_131) );
AO22x2_ASAP7_75t_L g132 ( .A1(n_102), .A2(n_84), .B1(n_85), .B2(n_88), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_102), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_119), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_102), .B(n_87), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_120), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_120), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_102), .B(n_79), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_108), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g143 ( .A(n_103), .B(n_74), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_99), .B(n_97), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_111), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_132), .A2(n_103), .B1(n_117), .B2(n_105), .Y(n_149) );
NOR2xp33_ASAP7_75t_R g150 ( .A(n_142), .B(n_111), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_127), .B(n_99), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_131), .B(n_104), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_144), .B(n_122), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_122), .B(n_116), .Y(n_154) );
NOR3xp33_ASAP7_75t_SL g155 ( .A(n_146), .B(n_114), .C(n_115), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_132), .A2(n_103), .B1(n_117), .B2(n_110), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_144), .B(n_101), .Y(n_159) );
NOR3xp33_ASAP7_75t_SL g160 ( .A(n_124), .B(n_107), .C(n_106), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_147), .A2(n_121), .B(n_98), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_144), .B(n_104), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_144), .B(n_118), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_132), .A2(n_110), .B1(n_112), .B2(n_121), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_122), .B(n_101), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_130), .B(n_110), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_131), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_143), .A2(n_112), .B1(n_98), .B2(n_100), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_122), .B(n_140), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_130), .A2(n_84), .B1(n_110), .B2(n_95), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_133), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_125), .Y(n_176) );
INVx3_ASAP7_75t_SL g177 ( .A(n_136), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_159), .B(n_130), .Y(n_184) );
AO32x1_ASAP7_75t_L g185 ( .A1(n_165), .A2(n_80), .A3(n_93), .B1(n_73), .B2(n_90), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_172), .Y(n_186) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_153), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_159), .B(n_153), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_172), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_172), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_157), .A2(n_136), .B1(n_140), .B2(n_110), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_177), .B(n_133), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_150), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_153), .B(n_133), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_173), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_161), .A2(n_139), .B(n_137), .C(n_126), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_159), .B(n_133), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_159), .B(n_133), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_157), .B(n_129), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_156), .A2(n_140), .B1(n_136), .B2(n_147), .Y(n_211) );
BUFx8_ASAP7_75t_L g212 ( .A(n_180), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_170), .B(n_136), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g217 ( .A(n_196), .B(n_160), .C(n_166), .Y(n_217) );
NAND2xp33_ASAP7_75t_L g218 ( .A(n_195), .B(n_140), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_214), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_187), .A2(n_149), .B1(n_170), .B2(n_162), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_195), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_182), .B(n_174), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_184), .A2(n_176), .B1(n_178), .B2(n_164), .Y(n_224) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_205), .A2(n_181), .B(n_179), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_214), .A2(n_174), .B1(n_152), .B2(n_151), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_183), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_212), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_188), .B(n_167), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_184), .A2(n_178), .B1(n_168), .B2(n_152), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_168), .B1(n_100), .B2(n_72), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_200), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_189), .B(n_140), .Y(n_234) );
CKINVDCx6p67_ASAP7_75t_R g235 ( .A(n_206), .Y(n_235) );
OAI21x1_ASAP7_75t_SL g236 ( .A1(n_182), .A2(n_175), .B(n_179), .Y(n_236) );
INVx6_ASAP7_75t_L g237 ( .A(n_212), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_189), .B(n_168), .Y(n_238) );
NAND2xp33_ASAP7_75t_SL g239 ( .A(n_213), .B(n_128), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_194), .A2(n_168), .B1(n_72), .B2(n_95), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_232), .A2(n_213), .B1(n_196), .B2(n_211), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_226), .B(n_209), .Y(n_243) );
AOI21xp33_ASAP7_75t_L g244 ( .A1(n_217), .A2(n_213), .B(n_211), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_223), .A2(n_205), .B(n_215), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_221), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_223), .A2(n_213), .B1(n_208), .B2(n_206), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_237), .A2(n_198), .B1(n_194), .B2(n_207), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_213), .B1(n_198), .B2(n_194), .Y(n_250) );
OAI211xp5_ASAP7_75t_L g251 ( .A1(n_219), .A2(n_155), .B(n_154), .C(n_86), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_237), .A2(n_208), .B1(n_206), .B2(n_193), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_193), .B1(n_190), .B2(n_188), .C(n_191), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_220), .A2(n_188), .B1(n_190), .B2(n_191), .C(n_186), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_227), .B(n_209), .Y(n_255) );
OAI322xp33_ASAP7_75t_L g256 ( .A1(n_240), .A2(n_86), .A3(n_75), .B1(n_97), .B2(n_192), .C1(n_197), .C2(n_210), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_237), .A2(n_207), .B1(n_198), .B2(n_168), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_188), .B1(n_190), .B2(n_186), .C(n_215), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_216), .B(n_209), .Y(n_261) );
AOI222xp33_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_75), .B1(n_210), .B2(n_197), .C1(n_192), .C2(n_207), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_235), .B(n_188), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_249), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_246), .B(n_238), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_243), .B(n_238), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_259), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_249), .B(n_238), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_262), .Y(n_269) );
AOI222xp33_ASAP7_75t_L g270 ( .A1(n_242), .A2(n_240), .B1(n_239), .B2(n_229), .C1(n_74), .C2(n_231), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_242), .A2(n_234), .B1(n_203), .B2(n_241), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_249), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_259), .A2(n_236), .B(n_179), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_246), .B(n_231), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_255), .B(n_239), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_248), .B(n_257), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_245), .B(n_241), .Y(n_278) );
NOR4xp25_ASAP7_75t_SL g279 ( .A(n_258), .B(n_90), .C(n_76), .D(n_78), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_245), .B(n_129), .Y(n_281) );
AOI322xp5_ASAP7_75t_L g282 ( .A1(n_255), .A2(n_233), .A3(n_137), .B1(n_139), .B2(n_82), .C1(n_79), .C2(n_73), .Y(n_282) );
AOI22xp33_ASAP7_75t_SL g283 ( .A1(n_250), .A2(n_212), .B1(n_233), .B2(n_218), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_260), .A2(n_165), .B(n_181), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_261), .B(n_229), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_267), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_278), .B(n_260), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_260), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_269), .A2(n_247), .B1(n_252), .B2(n_254), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
OAI211xp5_ASAP7_75t_SL g292 ( .A1(n_282), .A2(n_251), .B(n_262), .C(n_69), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_264), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_283), .B(n_249), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_278), .B(n_244), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_265), .B(n_249), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_265), .B(n_76), .Y(n_303) );
OAI33xp33_ASAP7_75t_L g304 ( .A1(n_269), .A2(n_80), .A3(n_93), .B1(n_89), .B2(n_82), .B3(n_78), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
OAI22xp5_ASAP7_75t_SL g306 ( .A1(n_283), .A2(n_253), .B1(n_263), .B2(n_256), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_89), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
OAI33xp33_ASAP7_75t_L g312 ( .A1(n_271), .A2(n_69), .A3(n_77), .B1(n_4), .B2(n_5), .B3(n_8), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_270), .A2(n_229), .B1(n_218), .B2(n_136), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_281), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_282), .B(n_138), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g316 ( .A1(n_271), .A2(n_208), .A3(n_206), .B(n_256), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_275), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_288), .B(n_266), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_306), .A2(n_270), .B1(n_277), .B2(n_266), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_303), .B(n_275), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_288), .B(n_266), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_317), .B(n_268), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_289), .B(n_275), .Y(n_323) );
AOI22x1_ASAP7_75t_L g324 ( .A1(n_296), .A2(n_268), .B1(n_77), .B2(n_272), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_268), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_299), .B(n_268), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_299), .B(n_268), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_303), .B(n_77), .C(n_279), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_301), .B(n_285), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_297), .B(n_285), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_285), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_305), .B(n_274), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_305), .B(n_274), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_310), .B(n_274), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_292), .B(n_2), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_309), .B(n_272), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_306), .Y(n_345) );
NAND2xp33_ASAP7_75t_SL g346 ( .A(n_309), .B(n_279), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_311), .B(n_3), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_311), .B(n_284), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_109), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_296), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_287), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_293), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_302), .B(n_109), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_290), .B(n_4), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_293), .B(n_5), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_298), .B(n_8), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_298), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_302), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_319), .A2(n_313), .B(n_295), .Y(n_363) );
NAND2xp33_ASAP7_75t_SL g364 ( .A(n_358), .B(n_298), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_357), .A2(n_312), .B1(n_304), .B2(n_315), .C1(n_300), .C2(n_307), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_362), .B(n_300), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_345), .A2(n_313), .B1(n_300), .B2(n_308), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_342), .B(n_327), .Y(n_368) );
OR2x6_ASAP7_75t_L g369 ( .A(n_334), .B(n_307), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_349), .A2(n_316), .B(n_308), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_334), .B(n_308), .Y(n_371) );
OAI322xp33_ASAP7_75t_L g372 ( .A1(n_333), .A2(n_316), .A3(n_10), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_323), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_323), .B(n_352), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_336), .B(n_9), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_341), .A2(n_138), .B1(n_190), .B2(n_204), .C(n_199), .Y(n_378) );
OAI21xp33_ASAP7_75t_L g379 ( .A1(n_334), .A2(n_128), .B(n_134), .Y(n_379) );
AOI22x1_ASAP7_75t_L g380 ( .A1(n_358), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_380) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_359), .A2(n_13), .A3(n_14), .B1(n_16), .B2(n_17), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_324), .A2(n_222), .B1(n_208), .B2(n_206), .Y(n_382) );
AOI31xp33_ASAP7_75t_L g383 ( .A1(n_346), .A2(n_185), .A3(n_18), .B(n_19), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_325), .B(n_17), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_335), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_318), .B(n_19), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_353), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_333), .A2(n_20), .A3(n_21), .B1(n_128), .B2(n_134), .C1(n_145), .C2(n_185), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_318), .B(n_20), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
OAI32xp33_ASAP7_75t_L g392 ( .A1(n_359), .A2(n_185), .A3(n_203), .B1(n_202), .B2(n_199), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_324), .A2(n_222), .B1(n_208), .B2(n_134), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_320), .A2(n_222), .B1(n_134), .B2(n_145), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_337), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_321), .B(n_145), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_326), .B(n_23), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_326), .B(n_26), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_321), .B(n_145), .Y(n_399) );
OAI21xp33_ASAP7_75t_SL g400 ( .A1(n_354), .A2(n_185), .B(n_203), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_331), .B(n_185), .C(n_212), .Y(n_401) );
OR2x6_ASAP7_75t_L g402 ( .A(n_344), .B(n_202), .Y(n_402) );
NAND2xp33_ASAP7_75t_L g403 ( .A(n_338), .B(n_136), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_329), .B(n_145), .Y(n_404) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_360), .B(n_31), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_322), .A2(n_136), .B1(n_140), .B2(n_212), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_353), .Y(n_407) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_338), .A2(n_185), .B1(n_203), .B2(n_201), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_322), .B1(n_329), .B2(n_325), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
INVx4_ASAP7_75t_SL g411 ( .A(n_369), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_363), .A2(n_322), .B1(n_339), .B2(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_375), .B(n_339), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_388), .B(n_340), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_395), .B(n_350), .Y(n_415) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_384), .B(n_355), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_403), .A2(n_360), .B(n_343), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_391), .B(n_355), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_366), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_373), .B(n_353), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_377), .B(n_350), .Y(n_421) );
XNOR2xp5_ASAP7_75t_L g422 ( .A(n_386), .B(n_351), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
NOR3xp33_ASAP7_75t_SL g424 ( .A(n_372), .B(n_361), .C(n_348), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_385), .B(n_361), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_407), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_365), .B(n_348), .Y(n_428) );
OAI221xp5_ASAP7_75t_SL g429 ( .A1(n_367), .A2(n_351), .B1(n_347), .B2(n_343), .C(n_356), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_387), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_396), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_404), .B(n_347), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_370), .B(n_356), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_383), .B(n_360), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_397), .B(n_332), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_381), .A2(n_332), .B1(n_330), .B2(n_201), .C(n_134), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_400), .B(n_330), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_371), .B(n_32), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_402), .Y(n_444) );
OAI322xp33_ASAP7_75t_L g445 ( .A1(n_398), .A2(n_134), .A3(n_145), .B1(n_185), .B2(n_181), .C1(n_165), .C2(n_190), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_410), .B(n_378), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_424), .A2(n_380), .B(n_401), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_419), .Y(n_448) );
NOR2x1p5_ASAP7_75t_L g449 ( .A(n_439), .B(n_371), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_402), .Y(n_450) );
NAND3x1_ASAP7_75t_L g451 ( .A(n_436), .B(n_406), .C(n_379), .Y(n_451) );
OA211x2_ASAP7_75t_L g452 ( .A1(n_436), .A2(n_405), .B(n_382), .C(n_400), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_428), .A2(n_393), .B1(n_394), .B2(n_389), .Y(n_453) );
OAI21xp33_ASAP7_75t_L g454 ( .A1(n_440), .A2(n_392), .B(n_204), .Y(n_454) );
CKINVDCx14_ASAP7_75t_R g455 ( .A(n_418), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_426), .A2(n_204), .B1(n_173), .B2(n_141), .C(n_135), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_444), .A2(n_202), .B1(n_204), .B2(n_195), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_412), .A2(n_173), .B1(n_175), .B2(n_195), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_416), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_435), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_424), .A2(n_141), .B(n_135), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_417), .A2(n_195), .B(n_173), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_423), .A2(n_33), .B1(n_40), .B2(n_43), .C1(n_45), .C2(n_46), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_446), .A2(n_441), .B1(n_409), .B2(n_423), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_457), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_447), .B(n_438), .C(n_429), .Y(n_470) );
NAND2xp33_ASAP7_75t_SL g471 ( .A(n_449), .B(n_442), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_460), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_464), .A2(n_429), .B(n_431), .C(n_443), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_463), .B(n_415), .Y(n_474) );
AOI22xp5_ASAP7_75t_SL g475 ( .A1(n_455), .A2(n_422), .B1(n_411), .B2(n_437), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_461), .B(n_462), .Y(n_476) );
NOR2xp33_ASAP7_75t_R g477 ( .A(n_448), .B(n_437), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_463), .B(n_415), .Y(n_478) );
NOR2xp33_ASAP7_75t_R g479 ( .A(n_450), .B(n_434), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_451), .A2(n_452), .B1(n_453), .B2(n_420), .Y(n_480) );
AOI211xp5_ASAP7_75t_L g481 ( .A1(n_454), .A2(n_432), .B(n_445), .C(n_433), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_465), .A2(n_427), .B(n_411), .C(n_50), .Y(n_482) );
XOR2xp5_ASAP7_75t_L g483 ( .A(n_459), .B(n_411), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_467), .B(n_56), .C(n_57), .D(n_58), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_458), .A2(n_456), .B(n_466), .Y(n_485) );
AOI211x1_ASAP7_75t_L g486 ( .A1(n_466), .A2(n_447), .B(n_440), .C(n_439), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_456), .A2(n_455), .B1(n_448), .B2(n_460), .Y(n_487) );
NAND4xp75_ASAP7_75t_L g488 ( .A(n_486), .B(n_480), .C(n_468), .D(n_475), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_487), .A2(n_470), .B1(n_471), .B2(n_473), .C(n_472), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_477), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_476), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_469), .B(n_474), .Y(n_492) );
AND4x1_ASAP7_75t_L g493 ( .A(n_490), .B(n_482), .C(n_481), .D(n_485), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_489), .A2(n_483), .B1(n_484), .B2(n_478), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_491), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_495), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_495), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_497), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_498), .A2(n_488), .B1(n_494), .B2(n_496), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_499), .A2(n_493), .B1(n_482), .B2(n_479), .C(n_492), .Y(n_500) );
endmodule