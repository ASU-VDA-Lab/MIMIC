module fake_jpeg_20244_n_324 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_0),
.CON(n_27),
.SN(n_27)
);

BUFx2_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_19),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_14),
.B1(n_21),
.B2(n_12),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_32),
.C(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_25),
.A2(n_14),
.B1(n_16),
.B2(n_12),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_36),
.B(n_40),
.C(n_34),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_58),
.B1(n_38),
.B2(n_57),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_28),
.B1(n_17),
.B2(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_58),
.B1(n_40),
.B2(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_40),
.B1(n_42),
.B2(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_82),
.B1(n_80),
.B2(n_62),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_0),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_45),
.B1(n_43),
.B2(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_36),
.C(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_77),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_35),
.C(n_37),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_58),
.B1(n_59),
.B2(n_37),
.Y(n_83)
);

OAI22x1_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_35),
.B1(n_44),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_43),
.B1(n_46),
.B2(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_50),
.B1(n_54),
.B2(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_0),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_32),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_0),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_31),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_102),
.B1(n_92),
.B2(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_105),
.B1(n_119),
.B2(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_64),
.B1(n_75),
.B2(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_67),
.C(n_75),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_19),
.C(n_33),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_70),
.B(n_68),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_91),
.B(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_68),
.B1(n_76),
.B2(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_68),
.B1(n_76),
.B2(n_30),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_95),
.B1(n_60),
.B2(n_61),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_18),
.B(n_11),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_83),
.A2(n_76),
.B1(n_81),
.B2(n_29),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_103),
.B1(n_60),
.B2(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_22),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_84),
.CI(n_94),
.CON(n_135),
.SN(n_135)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_96),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_84),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_154),
.C(n_159),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_96),
.B1(n_91),
.B2(n_90),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_165),
.Y(n_190)
);

OAI211xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_85),
.B(n_89),
.C(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_164),
.B1(n_166),
.B2(n_124),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_101),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_145),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_107),
.B1(n_112),
.B2(n_114),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_107),
.B1(n_130),
.B2(n_105),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_98),
.B(n_18),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_112),
.B(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_18),
.B(n_33),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_156),
.B(n_104),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_153),
.A2(n_157),
.B1(n_128),
.B2(n_131),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_18),
.B(n_11),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_19),
.C(n_20),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_20),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_119),
.C(n_105),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_0),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_1),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_153),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_159),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_128),
.B1(n_131),
.B2(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_123),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_188),
.B(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_122),
.C(n_110),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_186),
.C(n_196),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_193),
.B1(n_149),
.B2(n_158),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_110),
.B(n_130),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_137),
.B(n_126),
.CI(n_106),
.CON(n_183),
.SN(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_142),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_110),
.B1(n_119),
.B2(n_104),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_189),
.B1(n_191),
.B2(n_157),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_115),
.C(n_111),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_162),
.B1(n_163),
.B2(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_128),
.B1(n_2),
.B2(n_1),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_22),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_15),
.C(n_13),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_147),
.B(n_152),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_206),
.B1(n_170),
.B2(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_207),
.B1(n_193),
.B2(n_190),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_148),
.B(n_145),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_141),
.B1(n_138),
.B2(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_209),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_151),
.B1(n_132),
.B2(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_214),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_150),
.B(n_146),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_164),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_221),
.B1(n_167),
.B2(n_185),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_150),
.B(n_146),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_169),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_224),
.A2(n_228),
.B1(n_237),
.B2(n_213),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_169),
.C(n_186),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_234),
.C(n_238),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_195),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_225),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_132),
.B1(n_188),
.B2(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_177),
.C(n_167),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_180),
.B1(n_191),
.B2(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_183),
.C(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_187),
.B1(n_156),
.B2(n_134),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_228),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_197),
.CI(n_219),
.CON(n_245),
.SN(n_245)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_246),
.Y(n_276)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_254),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_262),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_252),
.A2(n_260),
.B1(n_261),
.B2(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_199),
.C(n_201),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_259),
.C(n_243),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_209),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_251),
.B1(n_254),
.B2(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_209),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_204),
.B(n_217),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_206),
.C(n_202),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_212),
.B1(n_198),
.B2(n_208),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_268),
.B1(n_261),
.B2(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_273),
.C(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_252),
.A2(n_236),
.B1(n_239),
.B2(n_222),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_239),
.B1(n_231),
.B2(n_232),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_243),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_203),
.C(n_15),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_203),
.C(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_1),
.C(n_2),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_6),
.C(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_245),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_260),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_2),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_273),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_4),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_291),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_269),
.B1(n_272),
.B2(n_265),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_6),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_265),
.C(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_290),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_6),
.B(n_7),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_8),
.B(n_9),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_278),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_285),
.B(n_280),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_10),
.B(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_6),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_307),
.B(n_312),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_8),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_8),
.B(n_9),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_311),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_8),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_304),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_315),
.B1(n_308),
.B2(n_300),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_297),
.C(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_10),
.C(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_10),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_10),
.Y(n_324)
);


endmodule