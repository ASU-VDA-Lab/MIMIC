module real_jpeg_33056_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_0),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_0),
.Y(n_375)
);

BUFx12f_ASAP7_75t_L g510 ( 
.A(n_0),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_62),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_1),
.B(n_141),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_1),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_1),
.B(n_276),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_1),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_1),
.B(n_373),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_3),
.B(n_303),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_3),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_3),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_3),
.B(n_323),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_3),
.B(n_461),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_3),
.B(n_373),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_247),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_4),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_4),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_4),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_4),
.B(n_72),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_4),
.B(n_464),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_5),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_8),
.Y(n_513)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_9),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g263 ( 
.A(n_10),
.B(n_264),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g307 ( 
.A(n_10),
.B(n_96),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_10),
.B(n_335),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_10),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_10),
.B(n_476),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_10),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_10),
.B(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_11),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_11),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_11),
.B(n_62),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_11),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_11),
.B(n_198),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_11),
.B(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_11),
.B(n_533),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_21),
.B(n_561),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_12),
.Y(n_563)
);

NAND2x1_ASAP7_75t_SL g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_13),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_13),
.B(n_98),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_14),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_68),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_15),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_16),
.Y(n_132)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_17),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_18),
.B(n_217),
.Y(n_216)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_18),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_18),
.B(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_18),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_18),
.B(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_18),
.B(n_481),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_18),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_18),
.B(n_508),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_19),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_19),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_19),
.B(n_212),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_19),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_19),
.B(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_175),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_174),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_145),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_25),
.B(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_107),
.C(n_122),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_26),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_75),
.B(n_106),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_27),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_46),
.C(n_59),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_28),
.B(n_46),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_29),
.B(n_35),
.C(n_39),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_33),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_43),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_44),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.C(n_53),
.Y(n_46)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_47),
.B(n_50),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_49),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_52),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_53),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_55),
.B(n_310),
.Y(n_457)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_57),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_58),
.Y(n_332)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_59),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_66),
.C(n_74),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_64),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_74),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_67),
.B1(n_110),
.B2(n_113),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_110),
.C(n_114),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_95),
.C(n_97),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_71),
.A2(n_74),
.B1(n_97),
.B2(n_215),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_73),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_73),
.Y(n_461)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_73),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_93),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_76),
.A2(n_77),
.B1(n_93),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2x1_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_82),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_88),
.C(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_86),
.Y(n_442)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_87),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_93),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.C(n_105),
.Y(n_93)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_95),
.Y(n_221)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_97),
.A2(n_211),
.B1(n_215),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_100),
.B(n_105),
.Y(n_190)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_102),
.Y(n_327)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_192),
.C(n_200),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_105),
.B(n_201),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_122),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_120),
.C(n_121),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_113),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_156),
.C(n_157),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_112),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_121),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_144),
.C(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_133),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_129),
.C(n_133),
.Y(n_147)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_143),
.B2(n_144),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_172),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_158),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_224),
.B(n_557),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_177),
.A2(n_559),
.B(n_560),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_222),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_178),
.B(n_222),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_185),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_183),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_191),
.C(n_206),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_191),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_192),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_193),
.B(n_194),
.Y(n_260)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_197),
.B(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_219),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_208),
.B(n_210),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_216),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_214),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_219),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_286),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_SL g559 ( 
.A(n_228),
.B(n_230),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_R g230 ( 
.A(n_231),
.B(n_234),
.C(n_237),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

XNOR2x2_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_238),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_261),
.C(n_283),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.C(n_259),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_244),
.C(n_259),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_244),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_252),
.B(n_257),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_249),
.B(n_258),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_252),
.Y(n_388)
);

INVx3_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_259),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_284),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_272),
.B(n_282),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.C(n_270),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_SL g340 ( 
.A(n_263),
.B(n_267),
.C(n_270),
.Y(n_340)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_270),
.B1(n_271),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_278),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_273),
.B(n_278),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_273),
.B(n_278),
.Y(n_341)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_277),
.Y(n_386)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_277),
.Y(n_482)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_396),
.B(n_554),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_348),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_288),
.A2(n_555),
.B(n_556),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_345),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_289),
.B(n_345),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.C(n_343),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_291),
.B(n_343),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_294),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_318),
.C(n_336),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_352),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.C(n_312),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_297),
.B(n_299),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_300),
.A2(n_301),
.B1(n_312),
.B2(n_313),
.Y(n_423)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_305),
.B(n_308),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_363),
.Y(n_362)
);

AOI21xp33_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_309),
.B(n_311),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_305),
.A2(n_306),
.B1(n_311),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_310),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OA21x2_ASAP7_75t_SL g407 ( 
.A1(n_313),
.A2(n_314),
.B(n_317),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_337),
.B1(n_338),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.C(n_333),
.Y(n_319)
);

XOR2x1_ASAP7_75t_L g392 ( 
.A(n_320),
.B(n_393),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.C(n_328),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_324),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_329),
.A2(n_330),
.B1(n_333),
.B2(n_334),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_394),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_349),
.B(n_394),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.C(n_359),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_355),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_387),
.C(n_390),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_360),
.A2(n_361),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.C(n_376),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_362),
.B(n_446),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_365),
.A2(n_376),
.B1(n_377),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_366),
.A2(n_367),
.B1(n_371),
.B2(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_375),
.Y(n_535)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_382),
.C(n_383),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_379),
.B1(n_383),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_382),
.B(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_391),
.B1(n_392),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_450),
.B(n_552),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_424),
.B(n_427),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_398),
.B(n_424),
.C(n_553),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_420),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_421),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.C(n_408),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_407),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_408),
.B(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_414),
.C(n_416),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_466),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_456)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_466)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_448),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_428),
.B(n_448),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_431),
.C(n_444),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_445),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.C(n_443),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_443),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.C(n_440),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_440),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_437),
.B(n_501),
.Y(n_500)
);

INVx3_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_442),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_469),
.B(n_551),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_467),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_452),
.B(n_467),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_465),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_453),
.B(n_549),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_465),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.C(n_458),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_457),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_495),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

AO22x1_ASAP7_75t_L g491 ( 
.A1(n_459),
.A2(n_460),
.B1(n_462),
.B2(n_463),
.Y(n_491)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_546),
.B(n_550),
.Y(n_469)
);

OAI21x1_ASAP7_75t_SL g470 ( 
.A1(n_471),
.A2(n_503),
.B(n_545),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_492),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_472),
.B(n_492),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_485),
.C(n_491),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_473),
.A2(n_474),
.B1(n_541),
.B2(n_543),
.Y(n_540)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_479),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_498),
.C(n_499),
.Y(n_497)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_485),
.A2(n_486),
.B1(n_491),
.B2(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_490),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_490),
.Y(n_521)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_491),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_496),
.B2(n_502),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_493),
.B(n_497),
.C(n_500),
.Y(n_547)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_496),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_538),
.B(n_544),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_522),
.B(n_537),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_514),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_506),
.B(n_514),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_511),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_511),
.Y(n_530)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx8_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_511),
.B(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_521),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_518),
.B2(n_520),
.Y(n_515)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_516),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_520),
.C(n_521),
.Y(n_539)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_531),
.B(n_536),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_530),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_530),
.Y(n_536)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx3_ASAP7_75t_SL g533 ( 
.A(n_534),
.Y(n_533)
);

INVx8_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_540),
.Y(n_544)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_541),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_548),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_564),
.Y(n_561)
);

CKINVDCx11_ASAP7_75t_R g562 ( 
.A(n_563),
.Y(n_562)
);


endmodule