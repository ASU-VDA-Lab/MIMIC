module fake_jpeg_22339_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_20;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_1),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_37),
.B1(n_26),
.B2(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_28),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_2),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_52),
.B1(n_56),
.B2(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_66),
.B1(n_70),
.B2(n_72),
.Y(n_97)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_37),
.B1(n_30),
.B2(n_29),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_37),
.B1(n_29),
.B2(n_35),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_75),
.B(n_54),
.Y(n_90)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_37),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_36),
.C(n_23),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_37),
.B1(n_29),
.B2(n_35),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_35),
.B1(n_17),
.B2(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_90),
.B1(n_34),
.B2(n_32),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_69),
.C(n_59),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_86),
.C(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_89),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_50),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_71),
.B(n_67),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_34),
.B1(n_42),
.B2(n_44),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_62),
.B1(n_64),
.B2(n_60),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_45),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_114),
.C(n_116),
.Y(n_124)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_74),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_92),
.B(n_97),
.Y(n_133)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_111),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_110),
.B1(n_77),
.B2(n_80),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_93),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_64),
.C(n_60),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_46),
.C(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_78),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_2),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_88),
.B(n_89),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_130),
.B(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_84),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_134),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_90),
.B(n_94),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_100),
.C(n_114),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_62),
.B1(n_17),
.B2(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_42),
.C(n_91),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

OAI31xp33_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_107),
.A3(n_102),
.B(n_92),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_125),
.B(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_119),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_92),
.CI(n_103),
.CON(n_145),
.SN(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_128),
.B1(n_119),
.B2(n_129),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_124),
.C(n_136),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_76),
.B1(n_17),
.B2(n_104),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_156),
.B1(n_157),
.B2(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_25),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_91),
.B1(n_104),
.B2(n_26),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_132),
.B1(n_138),
.B2(n_124),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_121),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_147),
.C(n_141),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_167),
.B(n_170),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_123),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_23),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_2),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_27),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_3),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_23),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_177),
.B(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_27),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_16),
.B1(n_22),
.B2(n_20),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_146),
.B1(n_151),
.B2(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_167),
.C(n_172),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_149),
.B1(n_140),
.B2(n_173),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_204),
.C(n_205),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_163),
.B1(n_145),
.B2(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_145),
.C(n_24),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_24),
.C(n_22),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_20),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_16),
.B(n_18),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_16),
.B(n_18),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_190),
.B(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_191),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_186),
.C(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_205),
.Y(n_225)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_216),
.C(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_225),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_229),
.B(n_4),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_198),
.B1(n_204),
.B2(n_189),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_181),
.C(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_4),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_223),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_181),
.B(n_15),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_217),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_215),
.A3(n_219),
.B1(n_15),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_232)
);

AOI31xp67_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_5),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_8),
.B(n_9),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_5),
.CI(n_6),
.CON(n_240),
.SN(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

OAI21x1_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_233),
.B(n_11),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_13),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_10),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_243),
.C(n_10),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_12),
.B1(n_217),
.B2(n_236),
.Y(n_249)
);


endmodule