module fake_jpeg_29028_n_506 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_506);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_506;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_9),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_70),
.Y(n_121)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_9),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_64),
.B(n_86),
.Y(n_155)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_76),
.Y(n_135)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_10),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_38),
.B(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_96),
.Y(n_159)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_25),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_8),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_32),
.Y(n_163)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_108),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_49),
.B1(n_31),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_136),
.B1(n_150),
.B2(n_60),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_25),
.B1(n_45),
.B2(n_43),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_123),
.A2(n_143),
.B1(n_147),
.B2(n_157),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_83),
.A2(n_42),
.B1(n_45),
.B2(n_43),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_128),
.A2(n_62),
.B1(n_58),
.B2(n_51),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_69),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_89),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_76),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_55),
.B(n_30),
.Y(n_168)
);

NOR2x1_ASAP7_75t_R g173 ( 
.A(n_163),
.B(n_55),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_179),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_98),
.B1(n_82),
.B2(n_84),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_174),
.A2(n_177),
.B1(n_186),
.B2(n_209),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_68),
.B1(n_54),
.B2(n_67),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_183),
.A2(n_160),
.B1(n_156),
.B2(n_148),
.Y(n_241)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_105),
.C(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_204),
.Y(n_242)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_191),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_161),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_199),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_128),
.A2(n_85),
.B1(n_92),
.B2(n_73),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_211),
.B1(n_157),
.B2(n_139),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_85),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_202),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_45),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_205),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_121),
.B(n_73),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_43),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_115),
.B(n_165),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_135),
.B(n_102),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_117),
.A2(n_35),
.B1(n_51),
.B2(n_4),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_129),
.A2(n_35),
.B1(n_51),
.B2(n_6),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_214),
.B1(n_221),
.B2(n_171),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_150),
.A2(n_35),
.B1(n_3),
.B2(n_6),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_137),
.B(n_12),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_222),
.Y(n_243)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx9p33_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_12),
.B1(n_3),
.B2(n_7),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_135),
.B(n_7),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_166),
.B1(n_118),
.B2(n_126),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_236),
.B1(n_249),
.B2(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_173),
.A2(n_126),
.B1(n_118),
.B2(n_148),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_238),
.A2(n_241),
.B(n_244),
.C(n_245),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_183),
.A2(n_134),
.B1(n_170),
.B2(n_169),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_183),
.A2(n_134),
.B1(n_149),
.B2(n_146),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_145),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_259),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_183),
.A2(n_145),
.B1(n_167),
.B2(n_144),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_217),
.A2(n_125),
.B1(n_7),
.B2(n_11),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_210),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_188),
.B(n_0),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_186),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_221),
.B1(n_191),
.B2(n_219),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_281),
.B1(n_284),
.B2(n_238),
.Y(n_308)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_251),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_267),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_269),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_177),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_271),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_181),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_227),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_283),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_194),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_279),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_187),
.C(n_172),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_247),
.C(n_229),
.Y(n_321)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_209),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_212),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_282),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_253),
.B(n_215),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_250),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_235),
.A2(n_198),
.B1(n_206),
.B2(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_193),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_239),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_SL g287 ( 
.A(n_242),
.B(n_211),
.C(n_192),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_245),
.B(n_244),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_176),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_257),
.B(n_250),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_249),
.A2(n_185),
.B(n_178),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_224),
.B(n_262),
.Y(n_315)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_180),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_233),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_311),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_271),
.B(n_253),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_301),
.B(n_266),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_288),
.B(n_279),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_257),
.B(n_241),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_310),
.B(n_283),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_236),
.C(n_223),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_308),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_225),
.B(n_241),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_264),
.B(n_247),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_286),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_315),
.A2(n_252),
.B(n_290),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_263),
.A2(n_228),
.B1(n_241),
.B2(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_232),
.B1(n_239),
.B2(n_237),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_291),
.A2(n_237),
.B1(n_203),
.B2(n_189),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_294),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_322),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_335),
.B(n_341),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_324),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_327),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_267),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_291),
.B1(n_268),
.B2(n_288),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_329),
.B1(n_297),
.B2(n_304),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_291),
.B1(n_289),
.B2(n_282),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_291),
.B(n_284),
.Y(n_330)
);

OAI21x1_ASAP7_75t_R g351 ( 
.A1(n_330),
.A2(n_323),
.B(n_338),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_293),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_349),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_299),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_295),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_273),
.C(n_276),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_336),
.B(n_331),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_312),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_302),
.A2(n_275),
.B(n_291),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_338),
.A2(n_345),
.B(n_346),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_281),
.B1(n_280),
.B2(n_270),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_339),
.A2(n_317),
.B1(n_307),
.B2(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_273),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_225),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_229),
.C(n_316),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_278),
.B(n_269),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_348),
.Y(n_363)
);

OAI211xp5_ASAP7_75t_L g349 ( 
.A1(n_298),
.A2(n_307),
.B(n_299),
.C(n_295),
.Y(n_349)
);

AO21x1_ASAP7_75t_SL g381 ( 
.A1(n_351),
.A2(n_373),
.B(n_348),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_372),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_301),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_355),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_357),
.A2(n_367),
.B1(n_369),
.B2(n_370),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_378),
.B(n_346),
.Y(n_390)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_297),
.B1(n_320),
.B2(n_319),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_330),
.B1(n_325),
.B2(n_335),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_326),
.A2(n_318),
.B1(n_296),
.B2(n_313),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_296),
.B1(n_313),
.B2(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_309),
.B(n_306),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_347),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_374),
.B(n_375),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_336),
.B(n_331),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_376),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_344),
.C(n_333),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_296),
.B(n_306),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_381),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_386),
.C(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_383),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_336),
.C(n_332),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_353),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_390),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_339),
.C(n_341),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_397),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_352),
.A2(n_337),
.B1(n_343),
.B2(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_230),
.Y(n_395)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_366),
.B(n_256),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_396),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_353),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_398),
.Y(n_406)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_399),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_362),
.B(n_256),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_400),
.A2(n_396),
.B(n_383),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_358),
.B(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_402),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_367),
.A2(n_274),
.B1(n_265),
.B2(n_234),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_350),
.B1(n_360),
.B2(n_365),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_274),
.B1(n_265),
.B2(n_260),
.Y(n_405)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_411),
.A2(n_421),
.B1(n_399),
.B2(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_377),
.C(n_354),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_424),
.C(n_427),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_380),
.A2(n_350),
.B1(n_351),
.B2(n_356),
.Y(n_421)
);

AOI21xp33_ASAP7_75t_L g423 ( 
.A1(n_394),
.A2(n_356),
.B(n_360),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_373),
.B(n_400),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_370),
.C(n_359),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_358),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_426),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_357),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_389),
.B(n_369),
.C(n_361),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_384),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_443),
.C(n_444),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_380),
.B1(n_388),
.B2(n_397),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_416),
.B1(n_409),
.B2(n_408),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_401),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_435),
.Y(n_450)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

XOR2x2_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_398),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_433),
.Y(n_447)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_419),
.B(n_391),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_439),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_392),
.B1(n_387),
.B2(n_385),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_390),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_411),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_385),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_381),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_379),
.C(n_387),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_403),
.B1(n_379),
.B2(n_373),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_445),
.A2(n_421),
.B1(n_414),
.B2(n_416),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_446),
.A2(n_452),
.B1(n_226),
.B2(n_231),
.Y(n_474)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_434),
.A2(n_414),
.B(n_408),
.Y(n_453)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_445),
.A2(n_415),
.B(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_406),
.C(n_415),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_461),
.C(n_436),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_440),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_433),
.A2(n_422),
.B(n_405),
.Y(n_460)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_226),
.C(n_260),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_459),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_468),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_449),
.A2(n_447),
.B1(n_456),
.B2(n_451),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_465),
.A2(n_475),
.B1(n_455),
.B2(n_457),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_443),
.Y(n_466)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_428),
.Y(n_467)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_448),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_431),
.B1(n_430),
.B2(n_260),
.Y(n_469)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_430),
.C(n_226),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_458),
.C(n_461),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_460),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_175),
.B1(n_230),
.B2(n_208),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_463),
.B(n_473),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_476),
.A2(n_464),
.B(n_466),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_484),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_478),
.A2(n_471),
.B(n_450),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_470),
.B(n_457),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_479),
.B(n_483),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_450),
.C(n_453),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_475),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_L g487 ( 
.A1(n_482),
.A2(n_464),
.B(n_455),
.Y(n_487)
);

OAI321xp33_ASAP7_75t_L g494 ( 
.A1(n_487),
.A2(n_493),
.A3(n_480),
.B1(n_484),
.B2(n_488),
.C(n_486),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_489),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_491),
.B(n_492),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_481),
.A2(n_474),
.B(n_465),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_208),
.C(n_231),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_493),
.B(n_483),
.C(n_485),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_495),
.C(n_248),
.Y(n_500)
);

AOI21xp33_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_231),
.B(n_248),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_499),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_500),
.C(n_248),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_182),
.C(n_197),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_503),
.A2(n_11),
.B(n_14),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_15),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_14),
.B(n_0),
.Y(n_506)
);


endmodule