module real_jpeg_23844_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_0),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_0),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_0),
.B(n_42),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_27),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_46),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_27),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_1),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_16),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_4),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_46),
.Y(n_61)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_9),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_9),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_46),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_9),
.B(n_27),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_9),
.B(n_42),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_11),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_91),
.Y(n_161)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_13),
.B(n_27),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_46),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_42),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_15),
.B(n_25),
.Y(n_169)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_108),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.C(n_40),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_23),
.B(n_122),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_23),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_26),
.CI(n_29),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_39),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_40),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_45),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_41),
.B(n_44),
.CI(n_45),
.CON(n_114),
.SN(n_114)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_46),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_93),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.C(n_82),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_80),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_111),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_83),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_83),
.B(n_187),
.C(n_190),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.CI(n_86),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_184)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_120),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.C(n_119),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_114),
.B(n_188),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_114),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_119),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_191),
.C(n_192),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_185),
.C(n_186),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_174),
.C(n_175),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_154),
.C(n_155),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_141),
.C(n_146),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_139),
.C(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_136),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_160),
.C(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_173),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);


endmodule