module fake_jpeg_29444_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_13),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_27),
.B1(n_14),
.B2(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_42),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_12),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_26),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_14),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_25),
.B1(n_1),
.B2(n_3),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_25),
.B1(n_17),
.B2(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_56),
.B1(n_75),
.B2(n_66),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_62),
.B(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_34),
.B(n_20),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_25),
.B1(n_17),
.B2(n_18),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_66),
.B1(n_77),
.B2(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_15),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_47),
.C(n_46),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_40),
.B1(n_31),
.B2(n_43),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_97),
.B1(n_52),
.B2(n_88),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_18),
.A3(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_98),
.B(n_103),
.C(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_15),
.B(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_101),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_0),
.B(n_9),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_10),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_11),
.CI(n_0),
.CON(n_103),
.SN(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_101),
.B1(n_98),
.B2(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_117),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_49),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_122),
.B(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_67),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_54),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_112),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_63),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_134),
.B1(n_68),
.B2(n_88),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_97),
.C(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_122),
.C(n_120),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_128),
.B(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_63),
.B1(n_68),
.B2(n_88),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_129),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_106),
.B(n_114),
.C(n_111),
.D(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_138),
.B(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_110),
.B(n_108),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_138),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_115),
.B(n_105),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_115),
.B1(n_122),
.B2(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_145),
.B1(n_134),
.B2(n_123),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_125),
.C(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.C(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_128),
.C(n_132),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_145),
.A2(n_142),
.B1(n_143),
.B2(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_160),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_141),
.B(n_140),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_147),
.B(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_133),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_164),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_149),
.B1(n_155),
.B2(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_165),
.B(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_116),
.A3(n_109),
.B1(n_113),
.B2(n_104),
.C1(n_121),
.C2(n_84),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_171),
.B(n_79),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_109),
.A3(n_104),
.B1(n_84),
.B2(n_81),
.C1(n_77),
.C2(n_59),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_81),
.C(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_102),
.Y(n_175)
);


endmodule