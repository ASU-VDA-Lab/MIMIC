module real_aes_3073_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_983, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_984, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_982, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_983;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_984;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_982;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_976;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_746;
wire n_532;
wire n_656;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_973;
wire n_504;
wire n_725;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_449;
wire n_754;
wire n_607;
wire n_417;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_598;
wire n_404;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_727;
wire n_649;
wire n_749;
wire n_385;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_831;
wire n_487;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_429;
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_0), .A2(n_163), .B1(n_620), .B2(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_1), .A2(n_127), .B1(n_421), .B2(n_551), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_2), .A2(n_200), .B1(n_459), .B2(n_460), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_3), .A2(n_306), .B1(n_709), .B2(n_715), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_4), .A2(n_16), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_5), .A2(n_116), .B1(n_409), .B2(n_414), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_6), .A2(n_102), .B1(n_459), .B2(n_460), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_7), .A2(n_329), .B1(n_830), .B2(n_831), .Y(n_829) );
AOI22xp5_ASAP7_75t_SL g885 ( .A1(n_8), .A2(n_358), .B1(n_699), .B2(n_760), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_9), .A2(n_292), .B1(n_511), .B2(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_10), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_11), .A2(n_68), .B1(n_506), .B2(n_768), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_12), .A2(n_88), .B1(n_496), .B2(n_697), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_13), .A2(n_167), .B1(n_465), .B2(n_676), .Y(n_862) );
AOI222xp33_ASAP7_75t_SL g656 ( .A1(n_14), .A2(n_38), .B1(n_144), .B2(n_530), .C1(n_657), .C2(n_658), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_15), .A2(n_308), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_17), .A2(n_126), .B1(n_421), .B2(n_425), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_18), .Y(n_874) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_19), .A2(n_164), .B1(n_184), .B2(n_381), .C1(n_399), .C2(n_403), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_20), .A2(n_170), .B1(n_409), .B2(n_496), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_21), .A2(n_218), .B1(n_475), .B2(n_476), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g570 ( .A1(n_22), .A2(n_115), .B1(n_269), .B2(n_463), .C1(n_571), .C2(n_573), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_23), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_24), .A2(n_74), .B1(n_466), .B2(n_588), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g589 ( .A1(n_25), .A2(n_327), .B1(n_353), .B2(n_421), .C1(n_571), .C2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_26), .A2(n_283), .B1(n_451), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_27), .A2(n_282), .B1(n_618), .B2(n_822), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_28), .A2(n_35), .B1(n_421), .B2(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_29), .B(n_751), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_30), .A2(n_91), .B1(n_174), .B2(n_465), .C1(n_572), .C2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_31), .A2(n_227), .B1(n_510), .B2(n_579), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_32), .A2(n_226), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_33), .A2(n_39), .B1(n_510), .B2(n_742), .Y(n_878) );
INVx1_ASAP7_75t_SL g388 ( .A(n_34), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_34), .B(n_42), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_36), .A2(n_141), .B1(n_409), .B2(n_496), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_37), .A2(n_92), .B1(n_421), .B2(n_491), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_40), .A2(n_355), .B1(n_478), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_41), .A2(n_252), .B1(n_539), .B2(n_540), .Y(n_538) );
AO22x2_ASAP7_75t_L g390 ( .A1(n_42), .A2(n_342), .B1(n_387), .B2(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_43), .B(n_751), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_44), .A2(n_242), .B1(n_443), .B2(n_446), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_45), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_46), .A2(n_270), .B1(n_421), .B2(n_425), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_47), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_48), .A2(n_206), .B1(n_449), .B2(n_452), .Y(n_901) );
OA22x2_ASAP7_75t_L g753 ( .A1(n_49), .A2(n_754), .B1(n_755), .B2(n_777), .Y(n_753) );
INVx1_ASAP7_75t_L g777 ( .A(n_49), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_50), .A2(n_349), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_51), .A2(n_232), .B1(n_610), .B2(n_697), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_52), .A2(n_81), .B1(n_496), .B2(n_635), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_53), .A2(n_272), .B1(n_510), .B2(n_579), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_54), .A2(n_339), .B1(n_502), .B2(n_768), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_55), .A2(n_273), .B1(n_605), .B2(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g389 ( .A(n_56), .Y(n_389) );
AO22x1_ASAP7_75t_L g513 ( .A1(n_57), .A2(n_162), .B1(n_514), .B2(n_516), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_58), .A2(n_224), .B1(n_449), .B2(n_451), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_59), .A2(n_238), .B1(n_536), .B2(n_672), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_60), .B(n_572), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_61), .A2(n_107), .B1(n_466), .B2(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_62), .A2(n_343), .B1(n_510), .B2(n_579), .Y(n_578) );
AOI222xp33_ASAP7_75t_L g965 ( .A1(n_63), .A2(n_207), .B1(n_233), .B2(n_599), .C1(n_607), .C2(n_966), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_64), .A2(n_230), .B1(n_437), .B2(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_65), .B(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_66), .A2(n_145), .B1(n_508), .B2(n_539), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_67), .A2(n_246), .B1(n_531), .B2(n_760), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_69), .A2(n_118), .B1(n_429), .B2(n_433), .Y(n_428) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_70), .A2(n_179), .B1(n_387), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_71), .A2(n_360), .B1(n_443), .B2(n_446), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_72), .A2(n_248), .B1(n_399), .B2(n_760), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_73), .A2(n_289), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_75), .A2(n_198), .B1(n_601), .B2(n_603), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_76), .A2(n_244), .B1(n_510), .B2(n_511), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_77), .A2(n_955), .B1(n_974), .B2(n_975), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_77), .Y(n_974) );
AOI222xp33_ASAP7_75t_L g950 ( .A1(n_78), .A2(n_951), .B1(n_969), .B2(n_973), .C1(n_976), .C2(n_979), .Y(n_950) );
XOR2xp5_ASAP7_75t_L g954 ( .A(n_78), .B(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_79), .A2(n_169), .B1(n_481), .B2(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_80), .B(n_381), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_82), .A2(n_130), .B1(n_449), .B2(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_83), .A2(n_133), .B1(n_435), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_84), .A2(n_239), .B1(n_472), .B2(n_473), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_85), .A2(n_274), .B1(n_767), .B2(n_768), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_86), .A2(n_331), .B1(n_540), .B2(n_542), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_87), .A2(n_356), .B1(n_548), .B2(n_590), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_89), .A2(n_155), .B1(n_414), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_90), .A2(n_123), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_93), .A2(n_333), .B1(n_481), .B2(n_482), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_94), .A2(n_199), .B1(n_547), .B2(n_605), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_95), .A2(n_278), .B1(n_551), .B2(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_96), .B(n_641), .Y(n_640) );
XOR2x2_ASAP7_75t_L g686 ( .A(n_97), .B(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_98), .A2(n_325), .B1(n_690), .B2(n_709), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_99), .A2(n_192), .B1(n_473), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_100), .A2(n_150), .B1(n_478), .B2(n_776), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_101), .B(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_103), .A2(n_241), .B1(n_506), .B2(n_508), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_104), .A2(n_260), .B1(n_462), .B2(n_679), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_105), .B(n_751), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_106), .A2(n_171), .B1(n_481), .B2(n_482), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_108), .A2(n_301), .B1(n_551), .B2(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_109), .A2(n_132), .B1(n_421), .B2(n_551), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_110), .A2(n_135), .B1(n_496), .B2(n_635), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_111), .A2(n_185), .B1(n_496), .B2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_112), .A2(n_202), .B1(n_429), .B2(n_540), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_113), .A2(n_323), .B1(n_503), .B2(n_535), .Y(n_924) );
AO22x2_ASAP7_75t_L g394 ( .A1(n_114), .A2(n_288), .B1(n_387), .B2(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_117), .A2(n_350), .B1(n_503), .B2(n_539), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_119), .A2(n_361), .B1(n_614), .B2(n_709), .Y(n_880) );
OA22x2_ASAP7_75t_L g556 ( .A1(n_120), .A2(n_557), .B1(n_558), .B2(n_574), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_120), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_121), .A2(n_219), .B1(n_435), .B2(n_506), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_122), .A2(n_245), .B1(n_510), .B2(n_742), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_124), .A2(n_258), .B1(n_690), .B2(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_125), .A2(n_256), .B1(n_437), .B2(n_776), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_128), .B(n_751), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_129), .A2(n_254), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_131), .A2(n_136), .B1(n_403), .B2(n_747), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_134), .A2(n_299), .B1(n_516), .B2(n_535), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_137), .A2(n_203), .B1(n_742), .B2(n_847), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_138), .A2(n_348), .B1(n_610), .B2(n_697), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_139), .A2(n_354), .B1(n_497), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_140), .A2(n_188), .B1(n_459), .B2(n_460), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_142), .A2(n_205), .B1(n_459), .B2(n_460), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_143), .A2(n_236), .B1(n_472), .B2(n_473), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_146), .A2(n_267), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_147), .A2(n_158), .B1(n_478), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_148), .A2(n_324), .B1(n_760), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_149), .A2(n_287), .B1(n_539), .B2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_151), .A2(n_275), .B1(n_542), .B2(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_152), .A2(n_263), .B1(n_825), .B2(n_826), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_153), .A2(n_320), .B1(n_475), .B2(n_476), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_154), .A2(n_319), .B1(n_830), .B2(n_845), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_156), .A2(n_201), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_157), .A2(n_211), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_159), .A2(n_212), .B1(n_543), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_160), .A2(n_229), .B1(n_446), .B2(n_510), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_161), .A2(n_341), .B1(n_465), .B2(n_466), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_165), .A2(n_210), .B1(n_462), .B2(n_679), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_166), .B(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_168), .A2(n_191), .B1(n_450), .B2(n_451), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_172), .A2(n_298), .B1(n_437), .B2(n_439), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_173), .A2(n_175), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_176), .A2(n_314), .B1(n_496), .B2(n_635), .Y(n_744) );
OA22x2_ASAP7_75t_L g453 ( .A1(n_177), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_177), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_178), .A2(n_318), .B1(n_439), .B2(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g938 ( .A(n_179), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_180), .A2(n_285), .B1(n_566), .B2(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_181), .A2(n_316), .B1(n_672), .B2(n_673), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_182), .A2(n_250), .B1(n_462), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_183), .A2(n_312), .B1(n_481), .B2(n_482), .Y(n_791) );
INVx1_ASAP7_75t_L g377 ( .A(n_186), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_187), .A2(n_366), .B1(n_443), .B2(n_564), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_189), .A2(n_284), .B1(n_763), .B2(n_764), .Y(n_762) );
OA22x2_ASAP7_75t_L g733 ( .A1(n_190), .A2(n_734), .B1(n_735), .B2(n_752), .Y(n_733) );
INVx1_ASAP7_75t_L g752 ( .A(n_190), .Y(n_752) );
INVx1_ASAP7_75t_L g639 ( .A(n_193), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_193), .A2(n_194), .B(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_193), .A2(n_652), .B1(n_660), .B2(n_984), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_194), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_195), .A2(n_265), .B1(n_446), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_196), .A2(n_243), .B1(n_503), .B2(n_692), .Y(n_691) );
OAI22x1_ASAP7_75t_SL g594 ( .A1(n_197), .A2(n_595), .B1(n_623), .B2(n_624), .Y(n_594) );
INVx1_ASAP7_75t_L g623 ( .A(n_197), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_204), .A2(n_213), .B1(n_510), .B2(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_208), .B(n_599), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_209), .A2(n_276), .B1(n_429), .B2(n_451), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_214), .A2(n_234), .B1(n_506), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g487 ( .A(n_215), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_216), .A2(n_300), .B1(n_621), .B2(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g948 ( .A(n_217), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_220), .A2(n_268), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_221), .A2(n_302), .B1(n_535), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_222), .A2(n_364), .B1(n_610), .B2(n_697), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_223), .A2(n_311), .B1(n_403), .B2(n_658), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_225), .A2(n_351), .B1(n_421), .B2(n_590), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_228), .A2(n_322), .B1(n_399), .B2(n_403), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_231), .A2(n_235), .B1(n_451), .B2(n_478), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_237), .A2(n_280), .B1(n_421), .B2(n_425), .Y(n_700) );
XNOR2x1_ASAP7_75t_L g894 ( .A(n_240), .B(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_247), .A2(n_303), .B1(n_672), .B2(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_249), .B(n_381), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_251), .A2(n_317), .B1(n_459), .B2(n_460), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_253), .A2(n_522), .B1(n_523), .B2(n_553), .Y(n_521) );
INVx1_ASAP7_75t_L g553 ( .A(n_253), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_255), .A2(n_363), .B1(n_526), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_257), .A2(n_330), .B1(n_760), .B2(n_800), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_259), .B(n_552), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_261), .A2(n_279), .B1(n_421), .B2(n_491), .Y(n_645) );
INVx1_ASAP7_75t_L g949 ( .A(n_262), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_264), .A2(n_332), .B1(n_616), .B2(n_618), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_266), .B(n_421), .Y(n_722) );
AO22x1_ASAP7_75t_L g795 ( .A1(n_271), .A2(n_796), .B1(n_809), .B2(n_810), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_271), .Y(n_809) );
XNOR2x1_ASAP7_75t_L g818 ( .A(n_277), .B(n_819), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_281), .A2(n_334), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_286), .A2(n_313), .B1(n_429), .B2(n_614), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_288), .B(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_290), .A2(n_328), .B1(n_443), .B2(n_564), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_291), .A2(n_362), .B1(n_529), .B2(n_747), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_293), .A2(n_337), .B1(n_449), .B2(n_508), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_294), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_295), .A2(n_344), .B1(n_497), .B2(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_296), .B(n_381), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_297), .A2(n_336), .B1(n_479), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_304), .A2(n_321), .B1(n_403), .B2(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
XNOR2x2_ASAP7_75t_L g782 ( .A(n_307), .B(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_309), .A2(n_326), .B1(n_475), .B2(n_476), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_310), .B(n_552), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_315), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_335), .A2(n_365), .B1(n_475), .B2(n_476), .Y(n_790) );
INVx1_ASAP7_75t_L g910 ( .A(n_338), .Y(n_910) );
XNOR2x1_ASAP7_75t_L g840 ( .A(n_340), .B(n_841), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_345), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_346), .A2(n_359), .B1(n_531), .B2(n_760), .Y(n_958) );
INVx1_ASAP7_75t_L g933 ( .A(n_347), .Y(n_933) );
NAND2xp5_ASAP7_75t_SL g947 ( .A(n_347), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g934 ( .A(n_352), .Y(n_934) );
AND2x2_ASAP7_75t_R g978 ( .A(n_352), .B(n_933), .Y(n_978) );
INVxp67_ASAP7_75t_L g946 ( .A(n_357), .Y(n_946) );
AOI21xp33_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_929), .B(n_940), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_814), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_SL g929 ( .A1(n_370), .A2(n_815), .B(n_930), .Y(n_929) );
XNOR2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_626), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_519), .B2(n_625), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_485), .B1(n_517), .B2(n_518), .Y(n_374) );
INVx2_ASAP7_75t_L g518 ( .A(n_375), .Y(n_518) );
AOI22x1_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_453), .B1(n_483), .B2(n_484), .Y(n_375) );
INVx1_ASAP7_75t_SL g484 ( .A(n_376), .Y(n_484) );
XNOR2x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_427), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_408), .C(n_420), .Y(n_379) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_381), .Y(n_758) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_SL g468 ( .A(n_382), .Y(n_468) );
INVx4_ASAP7_75t_SL g599 ( .A(n_382), .Y(n_599) );
INVx3_ASAP7_75t_L g657 ( .A(n_382), .Y(n_657) );
INVx4_ASAP7_75t_SL g751 ( .A(n_382), .Y(n_751) );
INVx6_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_392), .Y(n_383) );
AND2x4_ASAP7_75t_L g401 ( .A(n_384), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g410 ( .A(n_384), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g460 ( .A(n_384), .B(n_411), .Y(n_460) );
AND2x2_ASAP7_75t_L g466 ( .A(n_384), .B(n_402), .Y(n_466) );
AND2x4_ASAP7_75t_L g572 ( .A(n_384), .B(n_392), .Y(n_572) );
AND2x2_ASAP7_75t_L g676 ( .A(n_384), .B(n_402), .Y(n_676) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_390), .Y(n_384) );
INVx2_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
AND2x2_ASAP7_75t_L g418 ( .A(n_385), .B(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_385), .Y(n_424) );
OAI22x1_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_388), .B2(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g391 ( .A(n_387), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_387), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_387), .Y(n_398) );
AND2x2_ASAP7_75t_L g406 ( .A(n_390), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
BUFx2_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
AND2x4_ASAP7_75t_L g431 ( .A(n_392), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_392), .B(n_406), .Y(n_438) );
AND2x4_ASAP7_75t_L g450 ( .A(n_392), .B(n_418), .Y(n_450) );
AND2x6_ASAP7_75t_L g475 ( .A(n_392), .B(n_406), .Y(n_475) );
AND2x2_ASAP7_75t_L g481 ( .A(n_392), .B(n_418), .Y(n_481) );
AND2x2_ASAP7_75t_L g673 ( .A(n_392), .B(n_432), .Y(n_673) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g405 ( .A(n_394), .B(n_396), .Y(n_405) );
INVx1_ASAP7_75t_L g413 ( .A(n_394), .Y(n_413) );
AND2x2_ASAP7_75t_L g423 ( .A(n_394), .B(n_397), .Y(n_423) );
INVxp67_ASAP7_75t_L g402 ( .A(n_396), .Y(n_402) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_413), .Y(n_417) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g531 ( .A(n_400), .Y(n_531) );
INVx2_ASAP7_75t_L g603 ( .A(n_400), .Y(n_603) );
INVx2_ASAP7_75t_L g658 ( .A(n_400), .Y(n_658) );
INVx1_ASAP7_75t_L g699 ( .A(n_400), .Y(n_699) );
INVx2_ASAP7_75t_L g747 ( .A(n_400), .Y(n_747) );
INVx2_ASAP7_75t_L g800 ( .A(n_400), .Y(n_800) );
INVx6_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g602 ( .A(n_403), .Y(n_602) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_404), .Y(n_530) );
BUFx2_ASAP7_75t_L g746 ( .A(n_404), .Y(n_746) );
BUFx2_ASAP7_75t_L g760 ( .A(n_404), .Y(n_760) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g426 ( .A(n_405), .B(n_418), .Y(n_426) );
AND2x4_ASAP7_75t_L g435 ( .A(n_405), .B(n_432), .Y(n_435) );
AND2x4_ASAP7_75t_L g462 ( .A(n_405), .B(n_418), .Y(n_462) );
AND2x2_ASAP7_75t_L g465 ( .A(n_405), .B(n_406), .Y(n_465) );
AND2x2_ASAP7_75t_L g588 ( .A(n_405), .B(n_406), .Y(n_588) );
AND2x2_ASAP7_75t_L g672 ( .A(n_405), .B(n_432), .Y(n_672) );
AND2x2_ASAP7_75t_L g445 ( .A(n_406), .B(n_417), .Y(n_445) );
AND2x2_ASAP7_75t_L g472 ( .A(n_406), .B(n_417), .Y(n_472) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_406), .B(n_417), .Y(n_670) );
AND2x4_ASAP7_75t_L g432 ( .A(n_407), .B(n_419), .Y(n_432) );
BUFx2_ASAP7_75t_SL g764 ( .A(n_409), .Y(n_764) );
BUFx6f_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g498 ( .A(n_410), .Y(n_498) );
BUFx3_ASAP7_75t_L g635 ( .A(n_410), .Y(n_635) );
BUFx4f_ASAP7_75t_L g697 ( .A(n_410), .Y(n_697) );
INVx1_ASAP7_75t_L g889 ( .A(n_410), .Y(n_889) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g527 ( .A(n_415), .Y(n_527) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_416), .Y(n_496) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_416), .Y(n_610) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x4_ASAP7_75t_L g441 ( .A(n_417), .B(n_432), .Y(n_441) );
AND2x4_ASAP7_75t_L g459 ( .A(n_417), .B(n_418), .Y(n_459) );
AND2x6_ASAP7_75t_L g476 ( .A(n_417), .B(n_432), .Y(n_476) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g549 ( .A(n_422), .Y(n_549) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x4_ASAP7_75t_L g446 ( .A(n_423), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g452 ( .A(n_423), .B(n_432), .Y(n_452) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_423), .B(n_424), .Y(n_463) );
AND2x4_ASAP7_75t_L g473 ( .A(n_423), .B(n_447), .Y(n_473) );
AND2x4_ASAP7_75t_L g482 ( .A(n_423), .B(n_432), .Y(n_482) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_423), .B(n_424), .Y(n_679) );
BUFx5_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
BUFx3_ASAP7_75t_L g590 ( .A(n_426), .Y(n_590) );
BUFx3_ASAP7_75t_L g968 ( .A(n_426), .Y(n_968) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_436), .C(n_442), .D(n_448), .Y(n_427) );
BUFx2_ASAP7_75t_L g770 ( .A(n_429), .Y(n_770) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
INVx2_ASAP7_75t_SL g502 ( .A(n_430), .Y(n_502) );
INVx4_ASAP7_75t_L g536 ( .A(n_430), .Y(n_536) );
INVx3_ASAP7_75t_SL g581 ( .A(n_430), .Y(n_581) );
INVx2_ASAP7_75t_L g620 ( .A(n_430), .Y(n_620) );
INVx8_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g540 ( .A(n_434), .Y(n_540) );
INVx1_ASAP7_75t_L g739 ( .A(n_434), .Y(n_739) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
BUFx3_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_435), .Y(n_776) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_435), .Y(n_808) );
INVx2_ASAP7_75t_L g638 ( .A(n_437), .Y(n_638) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
BUFx2_ASAP7_75t_L g566 ( .A(n_438), .Y(n_566) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g516 ( .A(n_440), .Y(n_516) );
INVx2_ASAP7_75t_L g543 ( .A(n_440), .Y(n_543) );
INVx2_ASAP7_75t_L g614 ( .A(n_440), .Y(n_614) );
INVx2_ASAP7_75t_L g690 ( .A(n_440), .Y(n_690) );
INVx2_ASAP7_75t_SL g715 ( .A(n_440), .Y(n_715) );
INVx2_ASAP7_75t_L g831 ( .A(n_440), .Y(n_831) );
INVx1_ASAP7_75t_SL g845 ( .A(n_440), .Y(n_845) );
INVx8_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g617 ( .A(n_444), .Y(n_617) );
INVx2_ASAP7_75t_L g655 ( .A(n_444), .Y(n_655) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
BUFx3_ASAP7_75t_L g773 ( .A(n_445), .Y(n_773) );
INVx5_ASAP7_75t_SL g512 ( .A(n_446), .Y(n_512) );
BUFx3_ASAP7_75t_L g579 ( .A(n_446), .Y(n_579) );
BUFx2_ASAP7_75t_L g848 ( .A(n_446), .Y(n_848) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx6_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
BUFx3_ASAP7_75t_L g713 ( .A(n_450), .Y(n_713) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_451), .Y(n_621) );
BUFx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g504 ( .A(n_452), .Y(n_504) );
BUFx2_ASAP7_75t_SL g537 ( .A(n_452), .Y(n_537) );
BUFx2_ASAP7_75t_SL g826 ( .A(n_452), .Y(n_826) );
BUFx3_ASAP7_75t_L g882 ( .A(n_452), .Y(n_882) );
INVx3_ASAP7_75t_L g483 ( .A(n_453), .Y(n_483) );
AO22x2_ASAP7_75t_L g794 ( .A1(n_453), .A2(n_483), .B1(n_795), .B2(n_811), .Y(n_794) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_469), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .C(n_464), .D(n_467), .Y(n_457) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_462), .Y(n_573) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_468), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .C(n_480), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_479), .Y(n_828) );
INVx2_ASAP7_75t_L g517 ( .A(n_485), .Y(n_517) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
XNOR2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_489), .B(n_499), .Y(n_488) );
AND4x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .C(n_494), .D(n_495), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g551 ( .A(n_492), .Y(n_551) );
INVx2_ASAP7_75t_L g721 ( .A(n_492), .Y(n_721) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_496), .Y(n_763) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .C(n_509), .Y(n_500) );
BUFx2_ASAP7_75t_L g649 ( .A(n_502), .Y(n_649) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g768 ( .A(n_504), .Y(n_768) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g539 ( .A(n_507), .Y(n_539) );
INVx1_ASAP7_75t_SL g644 ( .A(n_507), .Y(n_644) );
INVx2_ASAP7_75t_L g692 ( .A(n_507), .Y(n_692) );
INVx2_ASAP7_75t_L g825 ( .A(n_507), .Y(n_825) );
BUFx2_ASAP7_75t_L g641 ( .A(n_508), .Y(n_641) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
INVx2_ASAP7_75t_L g618 ( .A(n_512), .Y(n_618) );
INVx3_ASAP7_75t_L g742 ( .A(n_512), .Y(n_742) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g542 ( .A(n_515), .Y(n_542) );
INVx2_ASAP7_75t_L g709 ( .A(n_515), .Y(n_709) );
INVx2_ASAP7_75t_SL g830 ( .A(n_515), .Y(n_830) );
INVx1_ASAP7_75t_L g625 ( .A(n_519), .Y(n_625) );
XNOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_554), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR3xp33_ASAP7_75t_SL g523 ( .A(n_524), .B(n_532), .C(n_544), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx4f_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
NAND4xp25_ASAP7_75t_SL g532 ( .A(n_533), .B(n_534), .C(n_538), .D(n_541), .Y(n_532) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_546), .B(n_550), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
INVx2_ASAP7_75t_L g749 ( .A(n_549), .Y(n_749) );
XNOR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_594), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_575), .B1(n_592), .B2(n_593), .Y(n_555) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
INVx2_ASAP7_75t_L g574 ( .A(n_558), .Y(n_574) );
NAND4xp75_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .C(n_567), .D(n_570), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
BUFx3_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g719 ( .A(n_572), .Y(n_719) );
INVx1_ASAP7_75t_SL g593 ( .A(n_575), .Y(n_593) );
XOR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_591), .Y(n_575) );
NAND4xp75_ASAP7_75t_L g576 ( .A(n_577), .B(n_582), .C(n_585), .D(n_589), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_590), .Y(n_605) );
INVx2_ASAP7_75t_SL g624 ( .A(n_595), .Y(n_624) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_611), .Y(n_595) );
NAND4xp25_ASAP7_75t_SL g596 ( .A(n_597), .B(n_600), .C(n_604), .D(n_608), .Y(n_596) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx6f_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_615), .C(n_619), .D(n_622), .Y(n_611) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
XOR2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_729), .Y(n_626) );
XOR2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_683), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_663), .B1(n_681), .B2(n_682), .Y(n_629) );
INVx2_ASAP7_75t_SL g681 ( .A(n_630), .Y(n_681) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_646), .Y(n_630) );
OAI222xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_639), .B1(n_640), .B2(n_642), .C1(n_982), .C2(n_983), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_632), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .Y(n_632) );
BUFx6f_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_640), .B(n_642), .C(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_643), .B(n_645), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B(n_659), .Y(n_646) );
INVx1_ASAP7_75t_L g662 ( .A(n_649), .Y(n_662) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g823 ( .A(n_655), .Y(n_823) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_655), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OA22x2_ASAP7_75t_L g702 ( .A1(n_663), .A2(n_664), .B1(n_703), .B2(n_704), .Y(n_702) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_L g682 ( .A(n_664), .Y(n_682) );
XNOR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_680), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_674), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .C(n_669), .D(n_671), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .C(n_678), .Y(n_674) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_702), .B1(n_727), .B2(n_728), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g728 ( .A(n_686), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g687 ( .A(n_688), .B(n_695), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .C(n_693), .D(n_694), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .C(n_700), .D(n_701), .Y(n_695) );
INVx2_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
XOR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_726), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_716), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_711), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_713), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_723), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_720), .C(n_722), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_780), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_753), .B1(n_778), .B2(n_779), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_732), .Y(n_779) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_743), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .C(n_740), .D(n_741), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .C(n_748), .D(n_750), .Y(n_743) );
INVx2_ASAP7_75t_L g778 ( .A(n_753), .Y(n_778) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_765), .Y(n_755) );
NAND4xp25_ASAP7_75t_SL g756 ( .A(n_757), .B(n_759), .C(n_761), .D(n_762), .Y(n_756) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .C(n_771), .D(n_774), .Y(n_765) );
BUFx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g915 ( .A(n_776), .Y(n_915) );
OA22x2_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_794), .B1(n_812), .B2(n_813), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g812 ( .A(n_782), .Y(n_812) );
OR2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_789), .Y(n_783) );
NAND4xp25_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .C(n_787), .D(n_788), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .C(n_792), .D(n_793), .Y(n_789) );
INVx1_ASAP7_75t_L g813 ( .A(n_794), .Y(n_813) );
INVx1_ASAP7_75t_SL g811 ( .A(n_795), .Y(n_811) );
INVx1_ASAP7_75t_SL g810 ( .A(n_796), .Y(n_810) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_803), .Y(n_796) );
NAND4xp25_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .C(n_801), .D(n_802), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .C(n_806), .D(n_807), .Y(n_803) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
XNOR2x1_ASAP7_75t_L g815 ( .A(n_816), .B(n_837), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_832), .Y(n_819) );
NAND4xp25_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_827), .D(n_829), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .C(n_835), .D(n_836), .Y(n_832) );
XNOR2x1_ASAP7_75t_L g837 ( .A(n_838), .B(n_892), .Y(n_837) );
AO22x2_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_855), .B2(n_856), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OR2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_850), .Y(n_841) );
NAND4xp25_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .C(n_846), .D(n_849), .Y(n_842) );
NAND4xp25_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .C(n_853), .D(n_854), .Y(n_850) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OA22x2_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_875), .B2(n_891), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
XOR2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_874), .Y(n_858) );
NAND2x1_ASAP7_75t_SL g859 ( .A(n_860), .B(n_867), .Y(n_859) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
NOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_871), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
INVx1_ASAP7_75t_SL g891 ( .A(n_875), .Y(n_891) );
XNOR2x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_890), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_883), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .C(n_880), .D(n_881), .Y(n_877) );
NAND4xp25_ASAP7_75t_SL g883 ( .A(n_884), .B(n_885), .C(n_886), .D(n_887), .Y(n_883) );
INVx2_ASAP7_75t_SL g888 ( .A(n_889), .Y(n_888) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_908), .B1(n_927), .B2(n_928), .Y(n_893) );
INVx2_ASAP7_75t_L g928 ( .A(n_894), .Y(n_928) );
NAND4xp75_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .C(n_902), .D(n_905), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
AND2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
AND2x2_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g927 ( .A(n_908), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_917), .B2(n_926), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
INVxp67_ASAP7_75t_SL g911 ( .A(n_912), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g926 ( .A(n_912), .B(n_918), .C(n_923), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_916), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OR2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_923), .Y(n_917) );
NAND4xp25_ASAP7_75t_SL g918 ( .A(n_919), .B(n_920), .C(n_921), .D(n_922), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
INVx2_ASAP7_75t_SL g930 ( .A(n_931), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_932), .B(n_935), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_932), .B(n_936), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g944 ( .A(n_934), .Y(n_944) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
OAI21xp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_949), .B(n_950), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_942), .Y(n_941) );
AND2x4_ASAP7_75t_SL g942 ( .A(n_943), .B(n_945), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
OR2x2_ASAP7_75t_L g980 ( .A(n_944), .B(n_945), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g975 ( .A(n_955), .Y(n_975) );
NAND4xp75_ASAP7_75t_SL g955 ( .A(n_956), .B(n_959), .C(n_962), .D(n_965), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .Y(n_956) );
AND2x2_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_964), .Y(n_962) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g969 ( .A(n_970), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_971), .Y(n_970) );
CKINVDCx6p67_ASAP7_75t_R g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_SL g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_980), .Y(n_979) );
endmodule