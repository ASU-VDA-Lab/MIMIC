module fake_jpeg_27389_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_33;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_29),
.B1(n_20),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_67),
.B1(n_53),
.B2(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_58),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_45),
.B1(n_44),
.B2(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_11),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_86),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_82),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_33),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_16),
.B(n_25),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_92),
.B(n_60),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_47),
.B1(n_42),
.B2(n_66),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_23),
.B1(n_16),
.B2(n_45),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_39),
.B(n_47),
.C(n_42),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_43),
.B1(n_35),
.B2(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_102),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_12),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_73),
.C(n_59),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_98),
.C(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_89),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_92),
.B1(n_89),
.B2(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_124),
.B1(n_95),
.B2(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_7),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_93),
.B1(n_84),
.B2(n_78),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_65),
.B(n_93),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_104),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_0),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_102),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_128),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_117),
.C(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_135),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_114),
.B(n_118),
.Y(n_147)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_82),
.B1(n_35),
.B2(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_145),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_122),
.B1(n_116),
.B2(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_4),
.B1(n_13),
.B2(n_14),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_136),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_136),
.Y(n_155)
);

AO221x1_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_82),
.B1(n_112),
.B2(n_4),
.C(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_131),
.B1(n_141),
.B2(n_129),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_155),
.A2(n_143),
.B(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_133),
.C(n_132),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_6),
.C(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_142),
.C(n_146),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_153),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_160),
.B(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_14),
.B(n_171),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_158),
.B1(n_148),
.B2(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_150),
.B(n_13),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);


endmodule