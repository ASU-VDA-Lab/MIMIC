module fake_aes_109_n_172 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_172, n_632);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_172;
output n_632;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_165;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g76 ( .A(n_11), .B(n_62), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_15), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_73), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_54), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_39), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_69), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_11), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_59), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_26), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_22), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_43), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_37), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_14), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_2), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_72), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_28), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_36), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_75), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_18), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_19), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_65), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_44), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_60), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_16), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_47), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_24), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_21), .B(n_68), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_66), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_23), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_78), .Y(n_122) );
NOR2xp33_ASAP7_75t_R g123 ( .A(n_109), .B(n_107), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_92), .B(n_0), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_82), .A2(n_34), .B(n_71), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_92), .B(n_0), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_107), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_121), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_79), .B(n_1), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_121), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
BUFx8_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_93), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_93), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_99), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_99), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_77), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_105), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_86), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_86), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_100), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_96), .B(n_1), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_123), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_125), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
UNKNOWN g172 ( );
INVx1_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
AO22x2_ASAP7_75t_L g177 ( .A1(n_124), .A2(n_105), .B1(n_112), .B2(n_111), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_157), .A2(n_97), .B1(n_98), .B2(n_114), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_161), .B(n_101), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_125), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_161), .B(n_80), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_137), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_124), .B(n_102), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_140), .B(n_76), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_144), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_126), .B(n_94), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_126), .B(n_116), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_156), .B(n_120), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_140), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_127), .A2(n_106), .B1(n_108), .B2(n_110), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_153), .B(n_81), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_145), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_125), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_127), .A2(n_119), .B(n_88), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_144), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_125), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
INVx5_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
BUFx6f_ASAP7_75t_SL g211 ( .A(n_144), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_131), .B(n_87), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_154), .B(n_117), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_128), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_128), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_184), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_192), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_192), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_166), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
NAND3xp33_ASAP7_75t_SL g224 ( .A(n_202), .B(n_159), .C(n_149), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_189), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_213), .B(n_129), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_213), .B(n_131), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_213), .B(n_138), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_189), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_213), .B(n_144), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_211), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_187), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_195), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_177), .A2(n_138), .B1(n_160), .B2(n_155), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_199), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_173), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_211), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_217), .Y(n_244) );
NOR2xp33_ASAP7_75t_R g245 ( .A(n_167), .B(n_148), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_185), .B(n_151), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_199), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_175), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_185), .B(n_151), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_217), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_194), .A2(n_152), .B(n_172), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_181), .B(n_139), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_191), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_177), .A2(n_160), .B1(n_155), .B2(n_143), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_185), .B(n_139), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_185), .B(n_162), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_203), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_211), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_204), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_179), .B(n_141), .C(n_143), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_191), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_186), .B(n_158), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_214), .B(n_150), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_200), .B(n_158), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_200), .B(n_2), .Y(n_272) );
NOR3xp33_ASAP7_75t_SL g273 ( .A(n_179), .B(n_3), .C(n_4), .Y(n_273) );
BUFx2_ASAP7_75t_SL g274 ( .A(n_176), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_178), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_177), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_265), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_220), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_277), .A2(n_177), .B1(n_194), .B2(n_206), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_223), .B(n_176), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_237), .A2(n_201), .B(n_197), .C(n_212), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_228), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_237), .A2(n_190), .B1(n_193), .B2(n_198), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_246), .B(n_183), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_246), .B(n_186), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_225), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_231), .A2(n_205), .B(n_182), .Y(n_291) );
CKINVDCx11_ASAP7_75t_R g292 ( .A(n_277), .Y(n_292) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_230), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_246), .B(n_186), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_246), .B(n_186), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_251), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_228), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_255), .B(n_217), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_228), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_251), .B(n_201), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_223), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_251), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_241), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_241), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_234), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_249), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_259), .A2(n_182), .B(n_170), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_251), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_233), .B(n_217), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_234), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_268), .B(n_197), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_270), .A2(n_205), .B(n_170), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_233), .B(n_176), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_239), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_250), .A2(n_205), .B(n_170), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_267), .B(n_212), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_250), .A2(n_205), .B(n_170), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_233), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_256), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_239), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_284), .A2(n_254), .B1(n_226), .B2(n_258), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_323), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_323), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_278), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_288), .B(n_267), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_318), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_317), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_290), .B(n_276), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_278), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_323), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_280), .A2(n_257), .B1(n_256), .B2(n_271), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_318), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
BUFx4f_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_325), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_294), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_293), .A2(n_257), .B1(n_218), .B2(n_262), .Y(n_342) );
AOI221x1_ASAP7_75t_L g343 ( .A1(n_316), .A2(n_170), .B1(n_182), .B2(n_205), .C(n_208), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_299), .A2(n_226), .B1(n_229), .B2(n_227), .Y(n_344) );
AOI21xp33_ASAP7_75t_L g345 ( .A1(n_314), .A2(n_218), .B(n_272), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_293), .Y(n_346) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_291), .B(n_264), .C(n_273), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_292), .Y(n_348) );
AOI332xp33_ASAP7_75t_L g349 ( .A1(n_281), .A2(n_266), .A3(n_226), .B1(n_229), .B2(n_227), .B3(n_216), .C1(n_215), .C2(n_275), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_280), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_299), .A2(n_227), .B1(n_229), .B2(n_275), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_315), .B(n_227), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_305), .A2(n_226), .B1(n_229), .B2(n_224), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_305), .A2(n_266), .B1(n_244), .B2(n_252), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_287), .B1(n_288), .B2(n_297), .C(n_289), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
OAI332xp33_ASAP7_75t_L g358 ( .A1(n_333), .A2(n_315), .A3(n_301), .B1(n_296), .B2(n_321), .B3(n_215), .C1(n_216), .C2(n_188), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_347), .A2(n_319), .B1(n_324), .B2(n_310), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_345), .A2(n_266), .B1(n_245), .B2(n_303), .C(n_301), .Y(n_360) );
INVx5_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_347), .B(n_285), .C(n_311), .Y(n_362) );
CKINVDCx11_ASAP7_75t_R g363 ( .A(n_346), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_353), .A2(n_312), .B1(n_309), .B2(n_298), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_342), .A2(n_310), .B1(n_324), .B2(n_319), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_336), .A2(n_322), .B(n_320), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_333), .A2(n_309), .B1(n_312), .B2(n_307), .C(n_303), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_353), .A2(n_307), .B1(n_282), .B2(n_279), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_329), .A2(n_266), .B1(n_271), .B2(n_282), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_313), .B1(n_244), .B2(n_252), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_354), .A2(n_313), .B1(n_244), .B2(n_252), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_330), .A2(n_313), .B1(n_279), .B2(n_233), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_352), .A2(n_313), .B1(n_243), .B2(n_300), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_336), .A2(n_304), .B(n_306), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_325), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_334), .A2(n_243), .B1(n_308), .B2(n_306), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_344), .A2(n_308), .B1(n_262), .B2(n_232), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_349), .A2(n_317), .B(n_300), .C(n_286), .Y(n_381) );
AOI21xp33_ASAP7_75t_SL g382 ( .A1(n_348), .A2(n_232), .B(n_5), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_365), .A2(n_339), .B1(n_332), .B2(n_338), .Y(n_384) );
NOR4xp25_ASAP7_75t_SL g385 ( .A(n_367), .B(n_349), .C(n_350), .D(n_351), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_372), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_356), .A2(n_351), .B1(n_350), .B2(n_339), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_369), .B(n_337), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_339), .B1(n_332), .B2(n_338), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_361), .B(n_337), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_340), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_378), .B(n_340), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_338), .B1(n_355), .B2(n_335), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_335), .B1(n_328), .B2(n_327), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_359), .A2(n_328), .B1(n_327), .B2(n_209), .C(n_180), .Y(n_396) );
NOR2x2_ASAP7_75t_L g397 ( .A(n_363), .B(n_174), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_359), .B(n_240), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_371), .B(n_240), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_362), .Y(n_401) );
INVx4_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_368), .B(n_371), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_374), .A2(n_188), .B1(n_174), .B2(n_180), .C(n_243), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_381), .B(n_248), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_358), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_377), .B(n_248), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_373), .A2(n_300), .B1(n_286), .B2(n_302), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_376), .A2(n_286), .B1(n_302), .B2(n_295), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_382), .B(n_343), .C(n_171), .D(n_169), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_375), .B(n_263), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_379), .A2(n_243), .B1(n_302), .B2(n_295), .Y(n_415) );
BUFx2_ASAP7_75t_SL g416 ( .A(n_402), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_410), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_401), .B(n_163), .C(n_164), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_4), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_386), .B(n_5), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_410), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_406), .A2(n_235), .B1(n_295), .B2(n_302), .C(n_263), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_410), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_410), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_393), .B(n_343), .Y(n_426) );
OAI33xp33_ASAP7_75t_L g427 ( .A1(n_389), .A2(n_163), .A3(n_164), .B1(n_168), .B2(n_169), .B3(n_171), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_393), .B(n_6), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_400), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_403), .B(n_7), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_401), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_388), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_403), .B(n_7), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_401), .B(n_8), .Y(n_436) );
OAI33xp33_ASAP7_75t_L g437 ( .A1(n_412), .A2(n_168), .A3(n_9), .B1(n_10), .B2(n_12), .B3(n_15), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_387), .A2(n_295), .B1(n_317), .B2(n_283), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_392), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_390), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
OAI31xp33_ASAP7_75t_SL g442 ( .A1(n_412), .A2(n_8), .A3(n_16), .B(n_269), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_390), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_414), .B(n_269), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_398), .B(n_261), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_402), .B(n_247), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_398), .B(n_261), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_407), .B(n_210), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
AOI211xp5_ASAP7_75t_L g455 ( .A1(n_387), .A2(n_235), .B(n_170), .C(n_182), .Y(n_455) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_397), .A2(n_260), .A3(n_253), .B(n_238), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_391), .B(n_408), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
INVx6_ASAP7_75t_L g459 ( .A(n_391), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_396), .A2(n_405), .B1(n_399), .B2(n_385), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_408), .B(n_260), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_457), .B(n_405), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_457), .B(n_399), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_432), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_457), .B(n_385), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_446), .B(n_395), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_442), .A2(n_384), .B(n_396), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_433), .B(n_394), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_418), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_444), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_434), .B(n_413), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_431), .A2(n_404), .B1(n_415), .B2(n_413), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_416), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_446), .B(n_411), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
OAI31xp33_ASAP7_75t_L g477 ( .A1(n_431), .A2(n_404), .A3(n_409), .B(n_235), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_456), .B(n_210), .C(n_182), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_444), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_461), .B(n_208), .Y(n_481) );
AND3x2_ASAP7_75t_L g482 ( .A(n_454), .B(n_253), .C(n_25), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_461), .B(n_208), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_450), .B(n_208), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_437), .A2(n_165), .B1(n_210), .B2(n_182), .C(n_205), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_435), .B(n_208), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_439), .B(n_210), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_450), .B(n_208), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_452), .B(n_20), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
NAND2xp33_ASAP7_75t_SL g493 ( .A(n_435), .B(n_247), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_453), .A2(n_235), .B(n_236), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_460), .A2(n_247), .B1(n_221), .B2(n_238), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_440), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_416), .B(n_274), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_440), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_422), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_455), .A2(n_247), .B(n_236), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_422), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_428), .B(n_165), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_424), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_420), .B(n_221), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_436), .A2(n_219), .B(n_165), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_452), .B(n_27), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_436), .A2(n_247), .B1(n_176), .B2(n_219), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_29), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_445), .B(n_274), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_420), .B(n_176), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_458), .B(n_31), .Y(n_514) );
NOR2xp33_ASAP7_75t_R g515 ( .A(n_459), .B(n_35), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_421), .B(n_176), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_498), .Y(n_517) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_474), .A2(n_421), .B(n_438), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_498), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_463), .B(n_459), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_497), .A2(n_459), .B1(n_426), .B2(n_451), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_464), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_471), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_471), .A2(n_459), .B1(n_449), .B2(n_430), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_490), .B(n_443), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_485), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_463), .B(n_443), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_512), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g530 ( .A1(n_482), .A2(n_451), .B(n_423), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_467), .A2(n_473), .B1(n_477), .B2(n_505), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_479), .B(n_430), .C(n_425), .Y(n_532) );
AOI322xp5_ASAP7_75t_L g533 ( .A1(n_467), .A2(n_425), .A3(n_424), .B1(n_427), .B2(n_165), .C1(n_451), .C2(n_48), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_485), .Y(n_534) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_493), .A2(n_419), .A3(n_40), .B(n_42), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_500), .B(n_38), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_497), .A2(n_45), .B(n_46), .Y(n_537) );
OAI211xp5_ASAP7_75t_SL g538 ( .A1(n_495), .A2(n_49), .B(n_50), .C(n_52), .Y(n_538) );
AOI22x1_ASAP7_75t_SL g539 ( .A1(n_480), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_497), .A2(n_58), .B1(n_63), .B2(n_64), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_500), .B(n_70), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_464), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_472), .B(n_74), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_497), .A2(n_480), .B1(n_511), .B2(n_478), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_466), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_470), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_466), .B(n_468), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_465), .B(n_462), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_465), .B(n_503), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_476), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_475), .Y(n_553) );
AOI21xp33_ASAP7_75t_L g554 ( .A1(n_503), .A2(n_488), .B(n_497), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_477), .B(n_484), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_491), .B(n_508), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_515), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_511), .A2(n_478), .B(n_486), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_491), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_508), .B(n_507), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_529), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_519), .Y(n_562) );
AOI222xp33_ASAP7_75t_L g563 ( .A1(n_531), .A2(n_506), .B1(n_494), .B2(n_513), .C1(n_516), .C2(n_510), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_531), .B(n_532), .C(n_527), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_547), .A2(n_509), .B1(n_514), .B2(n_510), .C(n_499), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_524), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_547), .B(n_484), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_553), .B(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_521), .B(n_499), .Y(n_569) );
OAI211xp5_ASAP7_75t_L g570 ( .A1(n_518), .A2(n_487), .B(n_514), .C(n_483), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_559), .B(n_492), .Y(n_571) );
NOR3xp33_ASAP7_75t_SL g572 ( .A(n_530), .B(n_501), .C(n_487), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_545), .B(n_489), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_528), .B(n_492), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_551), .B(n_481), .Y(n_575) );
NAND2xp33_ASAP7_75t_SL g576 ( .A(n_559), .B(n_483), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_552), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_517), .B(n_502), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_550), .B(n_502), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_550), .B(n_504), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_520), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_552), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_551), .B(n_504), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_548), .B(n_534), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_546), .Y(n_585) );
OR2x6_ASAP7_75t_L g586 ( .A(n_544), .B(n_522), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_526), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_523), .Y(n_588) );
NOR4xp25_ASAP7_75t_SL g589 ( .A(n_560), .B(n_554), .C(n_549), .D(n_539), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_587), .B(n_523), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_572), .A2(n_558), .B(n_560), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_581), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_569), .B(n_525), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_586), .A2(n_557), .B1(n_556), .B2(n_555), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_564), .B(n_533), .C(n_535), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_589), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_576), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_576), .A2(n_537), .B(n_540), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_561), .B(n_543), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
XNOR2xp5_ASAP7_75t_L g601 ( .A(n_580), .B(n_536), .Y(n_601) );
XOR2xp5_ASAP7_75t_L g602 ( .A(n_567), .B(n_541), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_586), .A2(n_538), .B1(n_542), .B2(n_571), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_579), .B(n_573), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_584), .A2(n_579), .B1(n_566), .B2(n_570), .C(n_583), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_586), .A2(n_571), .B1(n_572), .B2(n_578), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_592), .B(n_566), .Y(n_607) );
NOR2xp33_ASAP7_75t_R g608 ( .A(n_596), .B(n_584), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_590), .Y(n_609) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_606), .A2(n_591), .B(n_603), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_597), .A2(n_565), .B1(n_575), .B2(n_568), .Y(n_611) );
XOR2xp5_ASAP7_75t_L g612 ( .A(n_602), .B(n_574), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_596), .B(n_577), .Y(n_613) );
OAI211xp5_ASAP7_75t_SL g614 ( .A1(n_605), .A2(n_563), .B(n_585), .C(n_582), .Y(n_614) );
OAI211xp5_ASAP7_75t_L g615 ( .A1(n_594), .A2(n_577), .B(n_582), .C(n_588), .Y(n_615) );
AO22x1_ASAP7_75t_L g616 ( .A1(n_599), .A2(n_593), .B1(n_604), .B2(n_600), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_595), .A2(n_605), .B1(n_591), .B2(n_606), .C(n_596), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_599), .A2(n_601), .B(n_598), .Y(n_618) );
OAI211xp5_ASAP7_75t_SL g619 ( .A1(n_591), .A2(n_605), .B(n_594), .C(n_572), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_597), .A2(n_594), .B1(n_606), .B2(n_586), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_610), .B(n_613), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_617), .B(n_619), .C(n_620), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_618), .A2(n_611), .B1(n_615), .B2(n_614), .C(n_612), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_608), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_624), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_622), .B(n_609), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_621), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_625), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_626), .Y(n_629) );
NOR2xp67_ASAP7_75t_L g630 ( .A(n_628), .B(n_627), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_630), .A2(n_623), .B1(n_627), .B2(n_629), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_631), .A2(n_616), .B(n_607), .Y(n_632) );
endmodule