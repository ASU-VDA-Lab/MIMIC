module real_jpeg_29763_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_24),
.B1(n_30),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_1),
.A2(n_35),
.B1(n_39),
.B2(n_56),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_35),
.B1(n_39),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_22),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_4),
.A2(n_30),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_4),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_4),
.B(n_76),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_33),
.B1(n_125),
.B2(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_24),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_6),
.A2(n_35),
.B1(n_39),
.B2(n_49),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_24),
.B1(n_30),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_8),
.A2(n_35),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_35),
.B1(n_39),
.B2(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_24),
.B1(n_30),
.B2(n_53),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_9),
.A2(n_30),
.A3(n_39),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_22),
.B1(n_23),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_24),
.B1(n_30),
.B2(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_35),
.B1(n_39),
.B2(n_68),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_94),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_93),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_69),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_18),
.B(n_69),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.C(n_58),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_19),
.A2(n_20),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_32),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.A3(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_22),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_61),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_22),
.A2(n_23),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_62),
.Y(n_64)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_28),
.B(n_52),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_28),
.B(n_42),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_33),
.A2(n_37),
.B1(n_42),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_33),
.A2(n_42),
.B1(n_119),
.B2(n_125),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_34),
.A2(n_41),
.B1(n_44),
.B2(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_34),
.A2(n_41),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_35),
.B(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_35),
.B(n_131),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_46),
.A2(n_58),
.B1(n_59),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_52),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_52),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_85),
.B2(n_86),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_135),
.B(n_141),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_115),
.B(n_134),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_112),
.C(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_122),
.B(n_133),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_121),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_127),
.B(n_132),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);


endmodule