module fake_jpeg_8321_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_21),
.Y(n_29)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_19),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_22),
.B1(n_20),
.B2(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_17),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_24),
.B(n_21),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_36),
.C(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_35),
.B1(n_12),
.B2(n_15),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_12),
.B1(n_11),
.B2(n_16),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_10),
.C(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_R g41 ( 
.A(n_32),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_49),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_44),
.B(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_51),
.B1(n_16),
.B2(n_28),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_47),
.B(n_48),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_42),
.C(n_35),
.Y(n_60)
);

A2O1A1O1Ixp25_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_51),
.B(n_54),
.C(n_53),
.D(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_63),
.C(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_70),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_74),
.B(n_5),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_4),
.Y(n_77)
);


endmodule