module fake_jpeg_28018_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_61),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_30),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_60),
.Y(n_90)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_25),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_42),
.C(n_39),
.Y(n_87)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_30),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_28),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_27),
.B1(n_29),
.B2(n_37),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_109)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_38),
.B1(n_19),
.B2(n_18),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_38),
.B1(n_19),
.B2(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_38),
.B1(n_19),
.B2(n_44),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_42),
.CI(n_48),
.CON(n_120),
.SN(n_120)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_29),
.B1(n_27),
.B2(n_33),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_32),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_51),
.B1(n_46),
.B2(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_74),
.B1(n_51),
.B2(n_86),
.Y(n_142)
);

AO22x2_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_56),
.B1(n_42),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_57),
.B1(n_49),
.B2(n_80),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_82),
.B1(n_88),
.B2(n_86),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_65),
.C(n_66),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_66),
.C(n_56),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_20),
.Y(n_149)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_68),
.Y(n_128)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_86),
.B1(n_69),
.B2(n_85),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_90),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_141),
.B1(n_147),
.B2(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_94),
.B(n_91),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_24),
.B(n_26),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_75),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_100),
.B1(n_105),
.B2(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_143),
.B1(n_101),
.B2(n_104),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_153),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_84),
.CI(n_89),
.CON(n_145),
.SN(n_145)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_85),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_69),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_95),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_120),
.C(n_119),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_157),
.C(n_167),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_120),
.C(n_109),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_136),
.B1(n_138),
.B2(n_133),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_161),
.B1(n_171),
.B2(n_5),
.Y(n_214)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_173),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_131),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_176),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_116),
.C(n_115),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_104),
.B1(n_101),
.B2(n_53),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_172),
.B1(n_180),
.B2(n_34),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_182),
.B1(n_21),
.B2(n_4),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_33),
.B1(n_31),
.B2(n_17),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_43),
.B1(n_107),
.B2(n_26),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_107),
.C(n_42),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_21),
.C(n_4),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_127),
.B(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_34),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_31),
.B(n_32),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_184),
.B(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_26),
.B1(n_24),
.B2(n_42),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_124),
.A2(n_24),
.B1(n_31),
.B2(n_34),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_129),
.B(n_135),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_0),
.B(n_3),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_184),
.B(n_173),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_145),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_209),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_126),
.A3(n_140),
.B1(n_139),
.B2(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_198),
.B1(n_214),
.B2(n_154),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_0),
.B(n_4),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_210),
.B(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_204),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_200),
.B1(n_197),
.B2(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_164),
.C(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_182),
.B(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_10),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_10),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_157),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_163),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_0),
.B(n_5),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_5),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_175),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_217),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_161),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_218),
.A2(n_192),
.B(n_198),
.Y(n_253)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_239),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_223),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_154),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_228),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_186),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_168),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_234),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_168),
.B1(n_164),
.B2(n_163),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_199),
.B1(n_194),
.B2(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_211),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_195),
.B1(n_202),
.B2(n_205),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_210),
.B(n_191),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_253),
.B(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_252),
.B1(n_255),
.B2(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_201),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_258),
.B1(n_261),
.B2(n_222),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_160),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_227),
.C(n_216),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_221),
.C(n_234),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_232),
.C(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.C(n_271),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_228),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_191),
.C(n_213),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_241),
.C(n_236),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_242),
.B(n_229),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_250),
.B1(n_248),
.B2(n_242),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_256),
.CI(n_244),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_253),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_206),
.B(n_215),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_11),
.B(n_14),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_255),
.B1(n_257),
.B2(n_259),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_15),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_288),
.B1(n_289),
.B2(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_243),
.C(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_222),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_287),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_209),
.B1(n_12),
.B2(n_13),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_276),
.B1(n_272),
.B2(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_11),
.C(n_14),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_277),
.C(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_263),
.C(n_264),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_273),
.C(n_266),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_275),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_269),
.C(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_9),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_12),
.C(n_14),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_305),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_15),
.C(n_6),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_291),
.B1(n_281),
.B2(n_282),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_5),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_7),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_304),
.B1(n_6),
.B2(n_7),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_7),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_314),
.B(n_311),
.C(n_307),
.D(n_315),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_322),
.C(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_306),
.Y(n_329)
);


endmodule