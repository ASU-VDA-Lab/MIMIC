module real_jpeg_11256_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_58),
.B1(n_71),
.B2(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_71),
.B1(n_78),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_81),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_81),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_12),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_12),
.A2(n_56),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_12),
.B(n_82),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_12),
.A2(n_31),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_31),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_45),
.B1(n_95),
.B2(n_148),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_85),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_85),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_104),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_88),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_87),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_22),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_40),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_24),
.B(n_77),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_40),
.B1(n_138),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_24),
.A2(n_40),
.B1(n_161),
.B2(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_24),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_25),
.B(n_29),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_25),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_26),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_31),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_31),
.B(n_61),
.Y(n_178)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_32),
.A2(n_63),
.B1(n_173),
.B2(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_84),
.B(n_86),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_40),
.A2(n_171),
.B(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_41),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_45),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_45),
.A2(n_95),
.B1(n_130),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_45),
.A2(n_132),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_45),
.A2(n_48),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_46),
.B(n_49),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_46),
.A2(n_47),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_47),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.C(n_83),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_53),
.B1(n_83),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B1(n_65),
.B2(n_66),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_54),
.A2(n_59),
.B1(n_65),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_56),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_61),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g173 ( 
.A(n_56),
.B(n_77),
.CON(n_173),
.SN(n_173)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_66),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_60),
.A2(n_64),
.B1(n_115),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_77),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_75),
.B1(n_80),
.B2(n_99),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_72),
.B(n_77),
.C(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_84),
.B(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_95),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_105),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_204),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_108),
.Y(n_204)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_112),
.A2(n_113),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_200),
.B(n_205),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_183),
.B(n_199),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_166),
.B(n_182),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_155),
.B(n_165),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_144),
.B(n_154),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_133),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_143),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_143),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_153),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_167),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.CI(n_162),
.CON(n_158),
.SN(n_158)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_164),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_181),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_175),
.C(n_181),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_194),
.C(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);


endmodule