module fake_aes_7947_n_860 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_860);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_860;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_818;
wire n_844;
wire n_725;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g226 ( .A(n_116), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_83), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_199), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_24), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_28), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_28), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_109), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_181), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_61), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_206), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_145), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_209), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_124), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_117), .B(n_21), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_225), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_39), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_11), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_110), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_123), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_138), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_47), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_171), .B(n_157), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_148), .Y(n_252) );
BUFx10_ASAP7_75t_L g253 ( .A(n_136), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_203), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_127), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_169), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_214), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_95), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_113), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_118), .Y(n_261) );
XOR2xp5_ASAP7_75t_L g262 ( .A(n_147), .B(n_139), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_94), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_66), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_6), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_1), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_122), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_85), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_186), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_180), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_173), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_60), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_6), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_177), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_140), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_108), .B(n_193), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_151), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_217), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_41), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_0), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_159), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_29), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_67), .B(n_207), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_54), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_40), .Y(n_285) );
CKINVDCx14_ASAP7_75t_R g286 ( .A(n_56), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_38), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_125), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_115), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_137), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_189), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_119), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_144), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_129), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_188), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_101), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_156), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_223), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_194), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_34), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_211), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_20), .Y(n_302) );
BUFx8_ASAP7_75t_SL g303 ( .A(n_175), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_36), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_3), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_74), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_219), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_149), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_37), .Y(n_309) );
INVxp33_ASAP7_75t_SL g310 ( .A(n_17), .Y(n_310) );
CKINVDCx14_ASAP7_75t_R g311 ( .A(n_3), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_215), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_66), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_68), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_16), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_153), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_1), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_102), .B(n_114), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_56), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_102), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_30), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_205), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_33), .Y(n_323) );
CKINVDCx16_ASAP7_75t_R g324 ( .A(n_52), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_132), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_9), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_182), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_168), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_107), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_104), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_84), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_70), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_133), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_201), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_221), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_143), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_220), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_165), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_179), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_210), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_224), .Y(n_341) );
NOR2xp67_ASAP7_75t_L g342 ( .A(n_42), .B(n_126), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_146), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_97), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_226), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_226), .Y(n_346) );
OAI22x1_ASAP7_75t_SL g347 ( .A1(n_305), .A2(n_4), .B1(n_0), .B2(n_2), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_284), .B(n_5), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_229), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_286), .A2(n_8), .B1(n_5), .B2(n_7), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_264), .B(n_7), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_226), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_229), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_244), .Y(n_355) );
INVx5_ASAP7_75t_L g356 ( .A(n_226), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_242), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_253), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_242), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_244), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_247), .A2(n_106), .B(n_105), .Y(n_362) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_264), .B(n_9), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_311), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_249), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_253), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_253), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_261), .B(n_12), .Y(n_368) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_279), .B(n_13), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_279), .B(n_13), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_324), .A2(n_16), .B1(n_14), .B2(n_15), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_282), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_353), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_351), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_356), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_371), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_371), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_358), .B(n_228), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_371), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_370), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_371), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_358), .B(n_298), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_373), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_373), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_362), .A2(n_233), .B(n_232), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_366), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_345), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_366), .B(n_367), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_352), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_348), .A2(n_310), .B1(n_257), .B2(n_277), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_374), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_380), .B(n_367), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_386), .B(n_367), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_362), .B(n_369), .C(n_363), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_391), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_379), .B(n_236), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_386), .B(n_236), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g413 ( .A1(n_375), .A2(n_362), .B(n_239), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_377), .A2(n_363), .B1(n_369), .B2(n_368), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_394), .B(n_384), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_377), .B(n_260), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_400), .B(n_235), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_381), .B(n_349), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_349), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_378), .B(n_238), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_381), .B(n_354), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_383), .B(n_381), .Y(n_425) );
AND2x6_ASAP7_75t_SL g426 ( .A(n_400), .B(n_347), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_385), .A2(n_355), .B(n_361), .C(n_354), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_389), .B(n_254), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_376), .B(n_372), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_389), .B(n_355), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_376), .Y(n_431) );
BUFx5_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_390), .B(n_361), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_395), .B(n_365), .Y(n_436) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_388), .B(n_350), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_395), .B(n_227), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_392), .B(n_254), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_364), .B1(n_281), .B2(n_316), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_393), .B(n_234), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_396), .B(n_240), .Y(n_442) );
INVx8_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_398), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_398), .A2(n_230), .B1(n_245), .B2(n_231), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_399), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_401), .B(n_237), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_401), .B(n_274), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_401), .B(n_243), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_407), .B(n_372), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_413), .A2(n_248), .B(n_246), .Y(n_456) );
OR2x6_ASAP7_75t_SL g457 ( .A(n_426), .B(n_259), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_427), .A2(n_265), .B(n_266), .C(n_263), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_412), .B(n_277), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_406), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_405), .A2(n_252), .B(n_251), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_443), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_405), .A2(n_258), .B(n_256), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_419), .B(n_302), .C(n_285), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_418), .A2(n_271), .B(n_270), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_443), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_438), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_425), .A2(n_422), .B(n_430), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_421), .A2(n_291), .B(n_288), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_437), .B(n_320), .C(n_309), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_429), .B(n_331), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_429), .A2(n_331), .B1(n_262), .B2(n_330), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_404), .A2(n_332), .B1(n_323), .B2(n_268), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_417), .A2(n_272), .B(n_280), .C(n_273), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_435), .A2(n_293), .B(n_292), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
AO32x2_ASAP7_75t_L g483 ( .A1(n_431), .A2(n_342), .A3(n_241), .B1(n_357), .B2(n_346), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g485 ( .A1(n_411), .A2(n_318), .B(n_283), .C(n_269), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_423), .A2(n_295), .B(n_294), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_444), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_416), .A2(n_287), .B1(n_300), .B2(n_296), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_445), .B(n_306), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_446), .B(n_313), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_447), .A2(n_314), .B1(n_317), .B2(n_315), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_433), .Y(n_493) );
OA22x2_ASAP7_75t_L g494 ( .A1(n_434), .A2(n_442), .B1(n_441), .B2(n_321), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_432), .B(n_303), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_441), .B(n_326), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_443), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_451), .B(n_344), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_452), .B(n_267), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_453), .A2(n_319), .B(n_328), .C(n_327), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_450), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_448), .A2(n_333), .B(n_334), .C(n_329), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_428), .A2(n_336), .B1(n_337), .B2(n_335), .Y(n_504) );
INVx8_ASAP7_75t_L g505 ( .A(n_439), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_428), .A2(n_339), .B1(n_340), .B2(n_338), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_439), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_407), .B(n_325), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_413), .A2(n_343), .B(n_341), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_406), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_413), .A2(n_269), .B(n_247), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_403), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_439), .B(n_282), .Y(n_513) );
BUFx8_ASAP7_75t_L g514 ( .A(n_439), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_425), .A2(n_275), .B(n_307), .C(n_299), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_407), .B(n_278), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_428), .A2(n_282), .B1(n_290), .B2(n_289), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_439), .B(n_282), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_413), .A2(n_322), .B(n_307), .Y(n_519) );
OR2x6_ASAP7_75t_L g520 ( .A(n_439), .B(n_250), .Y(n_520) );
OAI22x1_ASAP7_75t_L g521 ( .A1(n_440), .A2(n_301), .B1(n_308), .B2(n_297), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_407), .B(n_312), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_512), .B(n_255), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_473), .A2(n_276), .B(n_255), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_477), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_504), .A2(n_506), .B1(n_490), .B2(n_484), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_494), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_462), .A2(n_357), .B(n_359), .C(n_346), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_465), .A2(n_360), .B(n_356), .Y(n_529) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_519), .A2(n_357), .A3(n_359), .B(n_360), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_456), .A2(n_509), .B(n_482), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_493), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_502), .A2(n_112), .B(n_111), .Y(n_533) );
AO31x2_ASAP7_75t_L g534 ( .A1(n_515), .A2(n_19), .A3(n_17), .B(n_18), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_463), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_463), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_500), .A2(n_459), .B(n_488), .C(n_503), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_487), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_472), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_478), .A2(n_21), .B1(n_19), .B2(n_20), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_476), .A2(n_25), .B1(n_22), .B2(n_23), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_513), .A2(n_26), .B(n_27), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_471), .A2(n_31), .B1(n_27), .B2(n_30), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_505), .Y(n_544) );
AOI211xp5_ASAP7_75t_L g545 ( .A1(n_466), .A2(n_33), .B(n_31), .C(n_32), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_454), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_546) );
AOI221x1_ASAP7_75t_L g547 ( .A1(n_517), .A2(n_521), .B1(n_481), .B2(n_498), .C(n_474), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_499), .A2(n_121), .B(n_120), .Y(n_548) );
AO31x2_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_45), .A3(n_43), .B(n_44), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_468), .B(n_44), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_485), .A2(n_47), .B(n_45), .C(n_46), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_507), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_489), .B(n_48), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_461), .Y(n_555) );
AOI31xp67_ASAP7_75t_L g556 ( .A1(n_470), .A2(n_130), .A3(n_131), .B(n_128), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_518), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_557) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_492), .A2(n_53), .A3(n_54), .B(n_55), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_475), .B(n_53), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_464), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_497), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_510), .A2(n_135), .B(n_134), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_514), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_460), .B(n_57), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_486), .A2(n_58), .B(n_59), .C(n_60), .Y(n_565) );
AOI21xp5_ASAP7_75t_SL g566 ( .A1(n_495), .A2(n_142), .B(n_141), .Y(n_566) );
AO31x2_ASAP7_75t_L g567 ( .A1(n_483), .A2(n_61), .A3(n_62), .B(n_63), .Y(n_567) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_497), .Y(n_568) );
AO32x1_ASAP7_75t_L g569 ( .A1(n_483), .A2(n_63), .A3(n_64), .B1(n_65), .B2(n_68), .Y(n_569) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_483), .A2(n_152), .B(n_150), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_508), .A2(n_65), .B(n_69), .C(n_71), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_479), .B(n_71), .Y(n_572) );
AO31x2_ASAP7_75t_L g573 ( .A1(n_469), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_573) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_501), .A2(n_167), .B(n_218), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_522), .A2(n_166), .B(n_216), .Y(n_575) );
AO31x2_ASAP7_75t_L g576 ( .A1(n_516), .A2(n_73), .A3(n_75), .B(n_76), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g577 ( .A1(n_520), .A2(n_76), .B(n_77), .C(n_78), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_458), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_458), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_457), .B(n_79), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_471), .Y(n_581) );
AO32x2_ASAP7_75t_L g582 ( .A1(n_517), .A2(n_79), .A3(n_80), .B1(n_81), .B2(n_82), .Y(n_582) );
BUFx10_ASAP7_75t_L g583 ( .A(n_463), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_480), .A2(n_80), .B(n_81), .C(n_83), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_493), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_473), .A2(n_172), .B(n_213), .Y(n_586) );
INVx8_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_511), .A2(n_170), .B(n_212), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_467), .A2(n_85), .B(n_86), .C(n_87), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_478), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_471), .B(n_89), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_477), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_477), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_455), .B(n_90), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_527), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_535), .B(n_90), .Y(n_596) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_547), .A2(n_91), .A3(n_92), .B(n_93), .Y(n_597) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_524), .A2(n_174), .B(n_208), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_551), .B(n_91), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_583), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_583), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_526), .B(n_93), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_586), .A2(n_164), .B(n_204), .Y(n_604) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_535), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_553), .B(n_96), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_555), .Y(n_607) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_552), .A2(n_98), .A3(n_99), .B(n_100), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_581), .B(n_98), .Y(n_609) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_528), .A2(n_99), .A3(n_100), .B(n_101), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_594), .B(n_103), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_587), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_574), .A2(n_178), .B(n_202), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_560), .Y(n_614) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_588), .A2(n_163), .B(n_200), .Y(n_615) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_580), .A2(n_154), .B(n_155), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_554), .B(n_161), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_532), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_585), .B(n_162), .Y(n_619) );
OAI21x1_ASAP7_75t_SL g620 ( .A1(n_542), .A2(n_183), .B(n_185), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_536), .B(n_187), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_563), .B(n_190), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_538), .B(n_525), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_592), .B(n_191), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_562), .A2(n_192), .B(n_195), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_591), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_593), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_549), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_539), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_544), .B(n_536), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_536), .Y(n_631) );
BUFx3_ASAP7_75t_L g632 ( .A(n_561), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_568), .Y(n_633) );
NOR2x1_ASAP7_75t_SL g634 ( .A(n_579), .B(n_557), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_549), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_549), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
AO31x2_ASAP7_75t_L g638 ( .A1(n_589), .A2(n_571), .A3(n_565), .B(n_575), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_558), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_558), .Y(n_640) );
AO31x2_ASAP7_75t_L g641 ( .A1(n_533), .A2(n_548), .A3(n_543), .B(n_564), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_534), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_578), .B(n_523), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_559), .B(n_572), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_567), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_576), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_529), .A2(n_546), .B(n_566), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_545), .B(n_541), .Y(n_648) );
AO31x2_ASAP7_75t_L g649 ( .A1(n_556), .A2(n_570), .A3(n_530), .B(n_569), .Y(n_649) );
OR2x6_ASAP7_75t_L g650 ( .A(n_577), .B(n_550), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_540), .B(n_590), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_573), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_576), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_573), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_573), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_576), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_582), .B(n_530), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_582), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_537), .A2(n_584), .B(n_551), .C(n_531), .Y(n_660) );
OR2x6_ASAP7_75t_L g661 ( .A(n_587), .B(n_505), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_526), .A2(n_506), .B1(n_504), .B2(n_428), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_527), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_527), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_527), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_531), .A2(n_473), .B(n_409), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_531), .A2(n_473), .B(n_409), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_633), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_603), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_607), .B(n_614), .Y(n_670) );
AOI21xp5_ASAP7_75t_SL g671 ( .A1(n_626), .A2(n_604), .B(n_634), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_603), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
INVx4_ASAP7_75t_L g674 ( .A(n_661), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_618), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_623), .Y(n_676) );
AO21x2_ASAP7_75t_L g677 ( .A1(n_628), .A2(n_636), .B(n_635), .Y(n_677) );
INVx5_ASAP7_75t_L g678 ( .A(n_661), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_644), .B(n_602), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_603), .B(n_605), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_649), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_606), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_599), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_637), .B(n_639), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_605), .Y(n_685) );
AOI21xp5_ASAP7_75t_SL g686 ( .A1(n_604), .A2(n_662), .B(n_609), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_605), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_640), .B(n_646), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_629), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_595), .Y(n_690) );
AO21x2_ASAP7_75t_L g691 ( .A1(n_666), .A2(n_667), .B(n_653), .Y(n_691) );
AO21x2_ASAP7_75t_L g692 ( .A1(n_667), .A2(n_656), .B(n_655), .Y(n_692) );
OR2x6_ASAP7_75t_L g693 ( .A(n_622), .B(n_650), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_663), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_664), .B(n_665), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_642), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_600), .Y(n_697) );
BUFx3_ASAP7_75t_L g698 ( .A(n_612), .Y(n_698) );
BUFx3_ASAP7_75t_L g699 ( .A(n_601), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_652), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_648), .A2(n_660), .B(n_651), .Y(n_701) );
AO21x2_ASAP7_75t_L g702 ( .A1(n_657), .A2(n_658), .B(n_659), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_654), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_645), .Y(n_704) );
INVx4_ASAP7_75t_L g705 ( .A(n_632), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_624), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_611), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_611), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_619), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_619), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_610), .Y(n_711) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_631), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_610), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_610), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_608), .B(n_597), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_608), .B(n_597), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_608), .B(n_597), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_630), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_643), .B(n_650), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_643), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_596), .Y(n_721) );
INVx4_ASAP7_75t_SL g722 ( .A(n_638), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_641), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_647), .B(n_598), .Y(n_724) );
INVx5_ASAP7_75t_L g725 ( .A(n_620), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_617), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_616), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_625), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_673), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_675), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_678), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_668), .B(n_598), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_690), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_694), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_719), .B(n_621), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_689), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_670), .Y(n_737) );
AND2x4_ASAP7_75t_L g738 ( .A(n_719), .B(n_613), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_679), .B(n_615), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_676), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_704), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_679), .B(n_715), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_688), .B(n_720), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_688), .B(n_684), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_715), .B(n_716), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_684), .B(n_701), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_716), .B(n_717), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_702), .B(n_691), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_685), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_695), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_717), .B(n_702), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_680), .Y(n_752) );
BUFx2_ASAP7_75t_L g753 ( .A(n_699), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_699), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_691), .B(n_707), .Y(n_755) );
OR2x2_ASAP7_75t_L g756 ( .A(n_708), .B(n_711), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_697), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_697), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_713), .B(n_714), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_674), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_677), .B(n_728), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_682), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_683), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_720), .B(n_722), .Y(n_764) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_700), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_722), .B(n_693), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_759), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_742), .B(n_723), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_729), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_742), .B(n_723), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_745), .B(n_723), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_755), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_745), .B(n_722), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_765), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_747), .B(n_692), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_733), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_734), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_756), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_751), .B(n_700), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_753), .Y(n_780) );
AND2x4_ASAP7_75t_L g781 ( .A(n_766), .B(n_724), .Y(n_781) );
AND2x4_ASAP7_75t_L g782 ( .A(n_766), .B(n_724), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_730), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_744), .B(n_696), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_764), .B(n_703), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_761), .B(n_743), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_743), .B(n_681), .Y(n_787) );
INVx5_ASAP7_75t_L g788 ( .A(n_731), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_750), .B(n_706), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_743), .B(n_681), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_754), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_737), .B(n_726), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_769), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_786), .B(n_736), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_776), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_772), .B(n_748), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_777), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_783), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_784), .B(n_746), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_767), .B(n_762), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_774), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_767), .B(n_763), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_791), .Y(n_803) );
INVx6_ASAP7_75t_L g804 ( .A(n_788), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_778), .B(n_740), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_780), .B(n_739), .Y(n_806) );
INVxp33_ASAP7_75t_L g807 ( .A(n_785), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_768), .B(n_739), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_768), .B(n_752), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_779), .B(n_741), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_770), .B(n_752), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_793), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_794), .B(n_771), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_795), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_797), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_798), .Y(n_816) );
INVx3_ASAP7_75t_L g817 ( .A(n_804), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_800), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_799), .B(n_775), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_800), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_802), .Y(n_821) );
OR2x6_ASAP7_75t_L g822 ( .A(n_804), .B(n_686), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_808), .B(n_806), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_802), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_805), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_809), .B(n_773), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_812), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_818), .B(n_796), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_823), .B(n_807), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_814), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_820), .B(n_796), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_815), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_816), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_821), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_824), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_825), .Y(n_836) );
INVx1_ASAP7_75t_SL g837 ( .A(n_817), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_828), .B(n_819), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_829), .B(n_813), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_831), .B(n_810), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_837), .A2(n_822), .B1(n_788), .B2(n_803), .Y(n_841) );
OAI211xp5_ASAP7_75t_SL g842 ( .A1(n_827), .A2(n_792), .B(n_671), .C(n_789), .Y(n_842) );
NOR3xp33_ASAP7_75t_L g843 ( .A(n_834), .B(n_727), .C(n_721), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_L g844 ( .A1(n_830), .A2(n_698), .B(n_758), .C(n_757), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_835), .A2(n_811), .B1(n_826), .B2(n_781), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_836), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_832), .A2(n_781), .B1(n_782), .B2(n_773), .Y(n_847) );
NAND3xp33_ASAP7_75t_SL g848 ( .A(n_833), .B(n_760), .C(n_801), .Y(n_848) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_842), .A2(n_848), .B1(n_847), .B2(n_845), .C(n_844), .Y(n_849) );
O2A1O1Ixp33_ASAP7_75t_L g850 ( .A1(n_841), .A2(n_846), .B(n_843), .C(n_838), .Y(n_850) );
NOR2xp67_ASAP7_75t_L g851 ( .A(n_840), .B(n_839), .Y(n_851) );
NOR3xp33_ASAP7_75t_L g852 ( .A(n_849), .B(n_705), .C(n_718), .Y(n_852) );
OAI21xp5_ASAP7_75t_L g853 ( .A1(n_852), .A2(n_850), .B(n_851), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g854 ( .A1(n_853), .A2(n_732), .B(n_735), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_854), .A2(n_709), .B(n_710), .Y(n_855) );
AOI21xp33_ASAP7_75t_L g856 ( .A1(n_855), .A2(n_669), .B(n_687), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_856), .A2(n_788), .B(n_725), .C(n_687), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_857), .A2(n_725), .B1(n_672), .B2(n_712), .C(n_749), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_858), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_859), .A2(n_738), .B1(n_790), .B2(n_787), .Y(n_860) );
endmodule