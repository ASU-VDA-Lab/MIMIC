module fake_netlist_1_11673_n_8 (n_3, n_1, n_2, n_0, n_8);
input n_3;
input n_1;
input n_2;
input n_0;
output n_8;
wire n_6;
wire n_4;
wire n_5;
wire n_7;
OAI22xp5_ASAP7_75t_L g4 ( .A1(n_1), .A2(n_0), .B1(n_3), .B2(n_2), .Y(n_4) );
OAI22xp5_ASAP7_75t_L g5 ( .A1(n_0), .A2(n_1), .B1(n_3), .B2(n_2), .Y(n_5) );
OR2x2_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
NAND4xp25_ASAP7_75t_SL g7 ( .A(n_6), .B(n_5), .C(n_1), .D(n_2), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
endmodule