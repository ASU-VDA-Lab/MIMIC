module fake_jpeg_30212_n_259 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_34),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_50),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_0),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_22),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_19),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_12),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_73),
.B1(n_87),
.B2(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_72),
.B(n_96),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_21),
.B1(n_25),
.B2(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_105),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_95),
.B1(n_31),
.B2(n_32),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_21),
.B1(n_25),
.B2(n_37),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_25),
.B1(n_37),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_37),
.B1(n_39),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_22),
.B1(n_30),
.B2(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_23),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_101),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_18),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_26),
.B(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_46),
.B1(n_56),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_75),
.B1(n_91),
.B2(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_111),
.Y(n_149)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_122),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_52),
.B1(n_43),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_85),
.B1(n_100),
.B2(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_31),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_66),
.B1(n_65),
.B2(n_48),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_112),
.A2(n_122),
.B1(n_114),
.B2(n_133),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_48),
.B1(n_63),
.B2(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_137),
.B1(n_84),
.B2(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_116),
.A2(n_127),
.B1(n_136),
.B2(n_134),
.Y(n_165)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_124),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_85),
.B1(n_79),
.B2(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_128),
.Y(n_140)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_8),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_138),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_11),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_12),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_112),
.Y(n_159)
);

FAx1_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_103),
.CI(n_91),
.CON(n_141),
.SN(n_141)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_139),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_147),
.B1(n_154),
.B2(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_157),
.B1(n_148),
.B2(n_141),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_92),
.B1(n_100),
.B2(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_141),
.B1(n_144),
.B2(n_142),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_102),
.C(n_104),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_156),
.C(n_125),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_78),
.B1(n_91),
.B2(n_112),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_126),
.B1(n_109),
.B2(n_130),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_123),
.B(n_111),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_162),
.B(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_117),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_121),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_169),
.B(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_171),
.Y(n_195)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_178),
.C(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_187),
.B1(n_189),
.B2(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_186),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_143),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_166),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_190),
.C(n_174),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_156),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_161),
.C(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_145),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_141),
.C(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_155),
.B1(n_151),
.B2(n_158),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_151),
.C(n_185),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_183),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_167),
.B(n_189),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_167),
.B(n_176),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_219),
.B(n_222),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_207),
.C(n_210),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_203),
.B1(n_169),
.B2(n_177),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_208),
.B(n_209),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_235),
.B(n_222),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_207),
.A3(n_200),
.B1(n_191),
.B2(n_197),
.C1(n_194),
.C2(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_188),
.B1(n_196),
.B2(n_169),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_216),
.B1(n_211),
.B2(n_217),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_196),
.B(n_193),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_233),
.B(n_231),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_223),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_195),
.Y(n_241)
);

AOI31xp67_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_223),
.A3(n_195),
.B(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_247),
.B(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_248),
.A2(n_225),
.B1(n_188),
.B2(n_192),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_231),
.B1(n_228),
.B2(n_238),
.Y(n_251)
);

AOI31xp67_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_237),
.A3(n_236),
.B(n_240),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_246),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_254),
.B(n_188),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_188),
.Y(n_259)
);


endmodule