module fake_jpeg_9369_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_0),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_40),
.B1(n_21),
.B2(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_25),
.B1(n_33),
.B2(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_37),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_41),
.B(n_24),
.C(n_34),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_26),
.CI(n_17),
.CON(n_124),
.SN(n_124)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_74),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_69),
.B1(n_68),
.B2(n_60),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_93),
.B1(n_69),
.B2(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_101),
.B1(n_62),
.B2(n_63),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_37),
.C(n_41),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_39),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_51),
.B1(n_31),
.B2(n_18),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_15),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_21),
.B1(n_24),
.B2(n_40),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_119),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_64),
.C(n_50),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_92),
.C(n_89),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_48),
.B1(n_68),
.B2(n_60),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_112),
.B1(n_51),
.B2(n_94),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_109),
.A2(n_75),
.B(n_99),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_36),
.A3(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_60),
.B1(n_51),
.B2(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_129),
.B1(n_76),
.B2(n_88),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_46),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_46),
.B(n_45),
.C(n_36),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_93),
.B1(n_84),
.B2(n_87),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_46),
.B(n_45),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_80),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_137),
.Y(n_167)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_130),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_139),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_142),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_152),
.Y(n_169)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_72),
.B1(n_94),
.B2(n_78),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_154),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_90),
.B1(n_95),
.B2(n_75),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_117),
.B1(n_122),
.B2(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_89),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_109),
.B(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_81),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_17),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_106),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_98),
.B1(n_86),
.B2(n_80),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_157),
.B1(n_163),
.B2(n_149),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_84),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_102),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_87),
.B1(n_85),
.B2(n_77),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_183),
.C(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_176),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_124),
.B(n_125),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_170),
.B(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_171),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_144),
.B1(n_162),
.B2(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_121),
.B(n_129),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_178),
.B(n_182),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_121),
.B1(n_126),
.B2(n_114),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_113),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_186),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_126),
.B1(n_110),
.B2(n_128),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_110),
.B(n_26),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_77),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_191),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_27),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_138),
.B1(n_132),
.B2(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_114),
.B1(n_115),
.B2(n_102),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_157),
.B1(n_140),
.B2(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_26),
.CI(n_85),
.CON(n_195),
.SN(n_195)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_26),
.Y(n_205)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_199),
.C(n_203),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_154),
.C(n_133),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_170),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_213),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_133),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_211),
.C(n_218),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_31),
.B1(n_133),
.B2(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_139),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_27),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_219),
.B(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_139),
.C(n_79),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_185),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_191),
.B1(n_188),
.B2(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_226),
.C(n_180),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_79),
.C(n_26),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_194),
.B1(n_176),
.B2(n_165),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_243),
.B1(n_210),
.B2(n_202),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_230),
.B(n_238),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_182),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_166),
.B1(n_177),
.B2(n_195),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_247),
.B1(n_249),
.B2(n_214),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_201),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_178),
.B1(n_195),
.B2(n_193),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_180),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_1),
.C(n_2),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_1),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_250),
.A2(n_216),
.B1(n_219),
.B2(n_202),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_27),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_27),
.C(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_210),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_224),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_257),
.B(n_227),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_208),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_218),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_214),
.B1(n_204),
.B2(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_204),
.B1(n_205),
.B2(n_226),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_268),
.B1(n_271),
.B2(n_235),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_269),
.B1(n_228),
.B2(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_27),
.Y(n_273)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

AOI211xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_229),
.B(n_238),
.C(n_252),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_283),
.B(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_254),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_289),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_237),
.B(n_245),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_270),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_273),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_258),
.C(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_250),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_298),
.C(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_250),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_296),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_270),
.B1(n_230),
.B2(n_264),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_267),
.C(n_261),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_272),
.B1(n_265),
.B2(n_251),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_6),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_8),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_290),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_6),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_305),
.B(n_275),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_274),
.B(n_279),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_284),
.A3(n_290),
.B1(n_286),
.B2(n_11),
.C(n_12),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_316),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_314),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_293),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_311),
.B(n_313),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_295),
.B1(n_10),
.B2(n_11),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_9),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_10),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_9),
.C(n_10),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_317),
.B1(n_10),
.B2(n_11),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_9),
.Y(n_326)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_12),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_332),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_12),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_323),
.C(n_322),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_330),
.B(n_318),
.C(n_331),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_333),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_328),
.B(n_13),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_13),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_14),
.C(n_271),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.Y(n_341)
);


endmodule