module real_jpeg_17917_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_576),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_0),
.B(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_1),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_2),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_49),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_49),
.B1(n_255),
.B2(n_259),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_3),
.A2(n_49),
.B1(n_276),
.B2(n_281),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_45),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_116),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_4),
.A2(n_116),
.B1(n_288),
.B2(n_292),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_4),
.A2(n_116),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_5),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_122),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_5),
.A2(n_122),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_5),
.A2(n_122),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_120),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_6),
.A2(n_191),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_6),
.A2(n_191),
.B1(n_255),
.B2(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_6),
.A2(n_191),
.B1(n_466),
.B2(n_469),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_7),
.Y(n_229)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_7),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_7),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_7),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_35),
.B1(n_81),
.B2(n_84),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_35),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_8),
.A2(n_35),
.B1(n_307),
.B2(n_310),
.Y(n_306)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_9),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_9),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_9),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_9),
.Y(n_445)
);

BUFx5_ASAP7_75t_L g500 ( 
.A(n_9),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_10),
.A2(n_166),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_10),
.A2(n_204),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_10),
.A2(n_204),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_10),
.A2(n_204),
.B1(n_494),
.B2(n_496),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_119),
.A3(n_207),
.B1(n_209),
.B2(n_215),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_12),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_12),
.A2(n_40),
.B1(n_214),
.B2(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_12),
.B(n_24),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_12),
.B(n_69),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_12),
.B(n_126),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_12),
.B(n_483),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_12),
.A2(n_210),
.B1(n_214),
.B2(n_267),
.Y(n_502)
);

OAI32xp33_ASAP7_75t_L g504 ( 
.A1(n_12),
.A2(n_505),
.A3(n_508),
.B1(n_511),
.B2(n_512),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_15),
.Y(n_577)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_16),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_16),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_16),
.Y(n_280)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_16),
.Y(n_481)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_155),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_153),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_22),
.B(n_62),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_23),
.A2(n_55),
.B(n_327),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OR2x6_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_44),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_24),
.A2(n_54),
.B1(n_187),
.B2(n_192),
.Y(n_186)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_26),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_27),
.Y(n_173)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_28),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_30),
.Y(n_507)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_34),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_42),
.Y(n_330)
);

OAI21x1_ASAP7_75t_SL g162 ( 
.A1(n_43),
.A2(n_112),
.B(n_117),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_48),
.Y(n_195)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_53),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_112),
.B1(n_117),
.B2(n_118),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_118),
.B(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_55),
.A2(n_117),
.B1(n_188),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_55),
.A2(n_117),
.B1(n_193),
.B2(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_55),
.A2(n_150),
.B(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_149),
.C(n_151),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_63),
.B(n_149),
.CI(n_151),
.CON(n_176),
.SN(n_176)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_110),
.C(n_124),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_64),
.A2(n_65),
.B1(n_124),
.B2(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_86),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_93),
.B(n_199),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_68),
.A2(n_94),
.B1(n_200),
.B2(n_266),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_68),
.A2(n_94),
.B1(n_266),
.B2(n_341),
.Y(n_340)
);

OAI22x1_ASAP7_75t_L g369 ( 
.A1(n_68),
.A2(n_94),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_68),
.A2(n_94),
.B1(n_341),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_95),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_69),
.A2(n_93),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_69),
.B(n_87),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_69),
.A2(n_93),
.B1(n_165),
.B2(n_390),
.Y(n_389)
);

AO22x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_73),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_137)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_75),
.Y(n_261)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_75),
.Y(n_291)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_80),
.A2(n_94),
.B(n_175),
.Y(n_331)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_87),
.Y(n_370)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_89),
.Y(n_343)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21x1_ASAP7_75t_SL g164 ( 
.A1(n_93),
.A2(n_165),
.B(n_174),
.Y(n_164)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_101),
.B2(n_106),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_109),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_114),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_162),
.C(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_125),
.B(n_164),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_136),
.B(n_144),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_126),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_126),
.B(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_126),
.A2(n_136),
.B1(n_421),
.B2(n_426),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_126),
.A2(n_136),
.B1(n_426),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_127),
.A2(n_251),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_127),
.B(n_145),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_127),
.A2(n_251),
.B1(n_492),
.B2(n_493),
.Y(n_491)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_131),
.B1(n_133),
.B2(n_135),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_129),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_133),
.Y(n_432)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_134),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_134),
.Y(n_457)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_134),
.Y(n_468)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_135),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_136),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_136),
.B(n_254),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_136),
.A2(n_392),
.B(n_534),
.Y(n_533)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_142),
.Y(n_428)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_143),
.Y(n_411)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_148),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_177),
.B(n_574),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_176),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_158),
.B(n_176),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_163),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_160),
.A2(n_162),
.B1(n_553),
.B2(n_554),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_160),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_162),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_162),
.A2(n_554),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_163),
.B(n_552),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_167),
.Y(n_372)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_173),
.Y(n_375)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g579 ( 
.A(n_176),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_549),
.B(n_571),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_543),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_401),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_355),
.C(n_381),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_333),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_297),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_183),
.B(n_297),
.C(n_545),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_249),
.C(n_270),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_184),
.B(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_205),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_198),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_186),
.B(n_198),
.C(n_205),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_196),
.A2(n_197),
.B1(n_442),
.B2(n_444),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_196),
.A2(n_197),
.B1(n_452),
.B2(n_456),
.Y(n_451)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_220),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_206),
.B(n_220),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_213),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_214),
.B(n_255),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_SL g421 ( 
.A1(n_214),
.A2(n_416),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_214),
.A2(n_222),
.B1(n_465),
.B2(n_472),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_214),
.B(n_408),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_230),
.B1(n_237),
.B2(n_242),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_221),
.A2(n_242),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_221),
.A2(n_450),
.B1(n_458),
.B2(n_459),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_221),
.A2(n_272),
.B(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_222),
.B(n_275),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_222),
.A2(n_306),
.B(n_362),
.Y(n_361)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_222),
.A2(n_431),
.B(n_438),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_222),
.A2(n_451),
.B1(n_465),
.B2(n_470),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_223),
.Y(n_469)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_225),
.Y(n_455)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_226),
.Y(n_362)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_229),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_230),
.A2(n_314),
.B(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_249),
.B(n_270),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_262),
.C(n_265),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_250),
.B(n_265),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_251),
.A2(n_253),
.B(n_317),
.Y(n_364)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_285),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_285),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_279),
.Y(n_437)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_296),
.Y(n_285)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_291),
.Y(n_510)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_322),
.C(n_332),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_322),
.B1(n_323),
.B2(n_332),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_315),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_301),
.B(n_315),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_314),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_302),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_306),
.Y(n_522)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_313),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_R g378 ( 
.A(n_324),
.B(n_326),
.C(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_353),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_334),
.B(n_353),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_339),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_335),
.B(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_339),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_346),
.C(n_348),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_340),
.B(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_348),
.Y(n_530)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g543 ( 
.A1(n_356),
.A2(n_544),
.B(n_546),
.C(n_547),
.D(n_548),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_357),
.B(n_358),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_377),
.B1(n_378),
.B2(n_380),
.Y(n_358)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_366),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_366),
.C(n_377),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_360)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_361),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_365),
.B1(n_397),
.B2(n_399),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_364),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g562 ( 
.A1(n_365),
.A2(n_399),
.B(n_563),
.Y(n_562)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_376),
.C(n_385),
.Y(n_384)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_376),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_381),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_382),
.B(n_383),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_384),
.B(n_387),
.C(n_395),
.Y(n_566)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_395),
.Y(n_386)
);

OA21x2_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_391),
.B(n_394),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_391),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_394),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_394),
.A2(n_557),
.B1(n_560),
.B2(n_570),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_397),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_400),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_537),
.B(n_542),
.Y(n_401)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_524),
.B(n_536),
.Y(n_402)
);

OAI21x1_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_487),
.B(n_523),
.Y(n_403)
);

AOI21x1_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_447),
.B(n_486),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_429),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_406),
.B(n_429),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_419),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_407),
.A2(n_419),
.B1(n_420),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_412),
.A3(n_414),
.B1(n_416),
.B2(n_417),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_418),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_439),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_440),
.C(n_446),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_446),
.Y(n_439)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_444),
.Y(n_495)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_462),
.B(n_485),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_460),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_460),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_475),
.B(n_484),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_474),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_474),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

BUFx12f_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_482),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_488),
.B(n_489),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_503),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_501),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_501),
.C(n_503),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_521),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_521),
.Y(n_532)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_SL g536 ( 
.A(n_525),
.B(n_526),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_531),
.B2(n_535),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_532),
.C(n_533),
.Y(n_541)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_531),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_541),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_565),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_550),
.A2(n_572),
.B(n_573),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_SL g550 ( 
.A(n_551),
.B(n_555),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_555),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_560),
.C(n_561),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_557),
.Y(n_570)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_558),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_561),
.A2(n_562),
.B1(n_568),
.B2(n_569),
.Y(n_567)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_SL g565 ( 
.A(n_566),
.B(n_567),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_566),
.B(n_567),
.Y(n_572)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);


endmodule