module real_jpeg_31761_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_714, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_714;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_704;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_703;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_712;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_699;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_708;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_0),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_0),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_2),
.A2(n_203),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_2),
.A2(n_203),
.B1(n_403),
.B2(n_407),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_2),
.A2(n_203),
.B1(n_510),
.B2(n_513),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_4),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_4),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_4),
.A2(n_291),
.B1(n_375),
.B2(n_377),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_4),
.A2(n_291),
.B1(n_480),
.B2(n_483),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_4),
.A2(n_291),
.B1(n_570),
.B2(n_573),
.Y(n_569)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_5),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_5),
.A2(n_143),
.B1(n_211),
.B2(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_5),
.A2(n_143),
.B1(n_276),
.B2(n_281),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_5),
.A2(n_143),
.B1(n_395),
.B2(n_397),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_6),
.A2(n_75),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_6),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_6),
.A2(n_342),
.B1(n_449),
.B2(n_453),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_6),
.A2(n_342),
.B1(n_541),
.B2(n_544),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_6),
.A2(n_342),
.B1(n_641),
.B2(n_643),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_7),
.A2(n_78),
.B1(n_130),
.B2(n_135),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_7),
.A2(n_78),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_7),
.A2(n_78),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_8),
.B(n_151),
.Y(n_426)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_8),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_8),
.B(n_70),
.Y(n_515)
);

OAI32xp33_ASAP7_75t_L g548 ( 
.A1(n_8),
.A2(n_549),
.A3(n_552),
.B1(n_554),
.B2(n_559),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_8),
.A2(n_476),
.B1(n_591),
.B2(n_594),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_L g622 ( 
.A1(n_8),
.A2(n_323),
.B(n_623),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_11),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_12),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_12),
.A2(n_150),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_12),
.A2(n_150),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_12),
.A2(n_150),
.B1(n_437),
.B2(n_440),
.Y(n_436)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_23),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_14),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_15),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_16),
.A2(n_385),
.B1(n_386),
.B2(n_389),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_16),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_16),
.A2(n_385),
.B1(n_490),
.B2(n_496),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_16),
.A2(n_385),
.B1(n_597),
.B2(n_599),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_16),
.A2(n_385),
.B1(n_611),
.B2(n_615),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_17),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_18),
.A2(n_59),
.B1(n_63),
.B2(n_67),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_18),
.A2(n_67),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_18),
.A2(n_67),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_708),
.Y(n_19)
);

AOI32xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_91),
.A3(n_354),
.B1(n_704),
.B2(n_705),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_22),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_22),
.B(n_712),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_24),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_89),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_87),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_27),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_27),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_27),
.B(n_95),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_57),
.B1(n_68),
.B2(n_71),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_29),
.A2(n_69),
.B(n_72),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_29),
.A2(n_69),
.B1(n_140),
.B2(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_29),
.A2(n_58),
.B1(n_69),
.B2(n_140),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_69),
.B1(n_146),
.B2(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2x1_ASAP7_75t_SL g288 ( 
.A(n_30),
.B(n_289),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_30),
.B(n_341),
.Y(n_340)
);

AO22x1_ASAP7_75t_L g383 ( 
.A1(n_30),
.A2(n_70),
.B1(n_341),
.B2(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_30),
.B(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_45),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_36),
.Y(n_422)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_37),
.Y(n_432)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_39),
.Y(n_345)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_40),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_40),
.Y(n_152)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_49),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_50),
.Y(n_159)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_50),
.Y(n_249)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_54),
.Y(n_429)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_56),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_56),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_62),
.Y(n_425)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_62),
.Y(n_475)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_67),
.A2(n_234),
.B(n_238),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_67),
.B(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_70),
.B(n_202),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_70),
.B(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_70),
.B(n_384),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_77),
.Y(n_390)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_84),
.Y(n_388)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_91),
.Y(n_710)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_221),
.C(n_300),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_191),
.Y(n_93)
);

AOI31xp33_ASAP7_75t_L g221 ( 
.A1(n_94),
.A2(n_222),
.A3(n_297),
.B(n_298),
.Y(n_221)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_94),
.B(n_297),
.C(n_301),
.D(n_353),
.Y(n_300)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_94),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_188),
.C(n_190),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_96),
.B(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_138),
.C(n_153),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_97),
.A2(n_98),
.B1(n_153),
.B2(n_154),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_97),
.A2(n_208),
.B(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_208),
.C(n_220),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_98),
.B(n_209),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_127),
.B(n_129),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_99),
.A2(n_127),
.B1(n_129),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_99),
.A2(n_479),
.B1(n_485),
.B2(n_486),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_99),
.B(n_673),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_99),
.A2(n_127),
.B1(n_479),
.B2(n_683),
.Y(n_682)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_100),
.A2(n_233),
.B1(n_275),
.B2(n_284),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_100),
.A2(n_275),
.B1(n_284),
.B2(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_100),
.A2(n_284),
.B1(n_308),
.B2(n_402),
.Y(n_401)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_100),
.A2(n_540),
.B(n_546),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_100),
.A2(n_284),
.B1(n_540),
.B2(n_596),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

OAI22x1_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_109),
.B2(n_112),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_103),
.Y(n_617)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_108),
.Y(n_658)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_110),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_112),
.Y(n_574)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_114),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_114),
.Y(n_572)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_114),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_115)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_116),
.Y(n_553)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_117),
.Y(n_484)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_123),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_123),
.Y(n_545)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_127),
.B(n_479),
.Y(n_546)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_128),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_128),
.B(n_476),
.Y(n_608)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_134),
.Y(n_311)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_134),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_134),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_149),
.Y(n_293)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_163),
.B1(n_179),
.B2(n_180),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_163),
.B1(n_210),
.B2(n_218),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_159),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_159),
.Y(n_331)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_159),
.Y(n_452)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_160),
.Y(n_181)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_179),
.B(n_180),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_163),
.A2(n_179),
.B1(n_210),
.B2(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_163),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_163),
.A2(n_218),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_163),
.B(n_521),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_167),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_172),
.B1(n_174),
.B2(n_178),
.Y(n_171)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_172),
.Y(n_453)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_179),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_179),
.B(n_374),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_179),
.B(n_489),
.Y(n_518)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_186),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_187),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_193),
.B(n_196),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_207),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_198),
.B(n_220),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_205),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_207),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g372 ( 
.A1(n_219),
.A2(n_328),
.B1(n_329),
.B2(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_219),
.B(n_476),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_295),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_223),
.B(n_295),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_294),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_225),
.B(n_230),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_251),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_230),
.A2(n_231),
.B(n_244),
.Y(n_352)
);

NAND2x1_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g598 ( 
.A(n_237),
.Y(n_598)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_242),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_243),
.Y(n_482)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_243),
.Y(n_664)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_248),
.Y(n_376)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

BUFx4f_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_269),
.B(n_285),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_252),
.A2(n_286),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_260),
.B(n_262),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_262),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_253),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_253),
.A2(n_326),
.B1(n_394),
.B2(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_253),
.B(n_569),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_253),
.A2(n_399),
.B1(n_638),
.B2(n_639),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

BUFx4f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_256),
.Y(n_396)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_256),
.Y(n_634)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_259),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_261),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_261),
.Y(n_628)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_267),
.Y(n_397)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_267),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_268),
.Y(n_439)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_268),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_268),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_269),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_270),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_271),
.Y(n_567)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_274),
.A2(n_350),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx4f_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_284),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_288),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_297),
.Y(n_702)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_302),
.B(n_304),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_R g304 ( 
.A(n_305),
.B(n_346),
.C(n_351),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_327),
.C(n_337),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_316),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_307),
.B(n_316),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_317),
.A2(n_323),
.B1(n_393),
.B2(n_398),
.Y(n_392)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_320),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22x1_ASAP7_75t_L g504 ( 
.A1(n_323),
.A2(n_436),
.B1(n_505),
.B2(n_509),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_323),
.A2(n_623),
.B(n_640),
.Y(n_680)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_337),
.B1(n_338),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_335),
.B2(n_336),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_328),
.A2(n_448),
.B(n_454),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_328),
.A2(n_454),
.B(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_339),
.B(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_352),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_353),
.B(n_701),
.Y(n_700)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_354),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_699),
.Y(n_354)
);

NAND2x1_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_529),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_455),
.B(n_525),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_358),
.B(n_696),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_361),
.B(n_408),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_359),
.B(n_361),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_359),
.B(n_361),
.Y(n_528)
);

MAJx2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.C(n_369),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_370),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_382),
.C(n_391),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_383),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_373),
.Y(n_521)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_378),
.Y(n_561)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_414),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_401),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_401),
.Y(n_466)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_400),
.Y(n_631)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_409),
.B(n_411),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_416),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_412),
.A2(n_413),
.B1(n_415),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_416),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_443),
.C(n_446),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_SL g462 ( 
.A(n_417),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_433),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_418),
.A2(n_419),
.B1(n_433),
.B2(n_434),
.Y(n_522)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

AOI32xp33_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.A3(n_423),
.B1(n_426),
.B2(n_427),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_441),
.Y(n_645)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_443),
.A2(n_444),
.B1(n_447),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_461),
.C(n_498),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g696 ( 
.A1(n_457),
.A2(n_697),
.B(n_698),
.Y(n_696)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_461),
.Y(n_697)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.C(n_467),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_466),
.B(n_468),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

MAJx2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_478),
.C(n_487),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_469),
.B(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_472),
.A2(n_476),
.B(n_477),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_476),
.B(n_555),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_476),
.B(n_631),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_476),
.B(n_661),
.Y(n_660)
);

OAI21xp33_ASAP7_75t_SL g673 ( 
.A1(n_476),
.A2(n_660),
.B(n_674),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_487),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_482),
.Y(n_603)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_523),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_499),
.B(n_523),
.Y(n_698)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.C(n_522),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_500),
.B(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_503),
.A2(n_522),
.B1(n_577),
.B2(n_578),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_515),
.B1(n_516),
.B2(n_519),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_515),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_515),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_504),
.A2(n_515),
.B1(n_516),
.B2(n_519),
.Y(n_579)
);

INVx3_ASAP7_75t_SL g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_509),
.A2(n_567),
.B(n_568),
.Y(n_566)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_520),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_522),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_527),
.B(n_528),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_695),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_580),
.B(n_693),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_575),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_533),
.B(n_694),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_538),
.C(n_547),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_583),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_537),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_538),
.A2(n_539),
.B1(n_547),
.B2(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_542),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_546),
.B(n_672),
.Y(n_671)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_566),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_566),
.Y(n_587)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_558),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_562),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_568),
.A2(n_610),
.B(n_618),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_575),
.Y(n_694)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_581),
.A2(n_604),
.B(n_692),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_582),
.B(n_585),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_582),
.B(n_585),
.Y(n_692)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_588),
.C(n_595),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_678),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g678 ( 
.A(n_589),
.B(n_595),
.Y(n_678)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_596),
.Y(n_683)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

OAI321xp33_ASAP7_75t_L g604 ( 
.A1(n_605),
.A2(n_676),
.A3(n_685),
.B1(n_690),
.B2(n_691),
.C(n_714),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_636),
.B(n_675),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_607),
.A2(n_621),
.B(n_635),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_609),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_608),
.B(n_609),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_610),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

BUFx2_ASAP7_75t_SL g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_622),
.B(n_629),
.Y(n_621)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_630),
.B(n_632),
.Y(n_629)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_637),
.B(n_646),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_637),
.B(n_646),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_647),
.B(n_671),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_647),
.B(n_671),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_648),
.A2(n_659),
.B1(n_665),
.B2(n_670),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_649),
.B(n_653),
.Y(n_648)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_649),
.Y(n_670)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

INVx6_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_666),
.B(n_668),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_667),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_669),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_677),
.B(n_679),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_677),
.B(n_679),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_680),
.B(n_681),
.C(n_684),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g687 ( 
.A(n_680),
.B(n_688),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_682),
.B1(n_684),
.B2(n_689),
.Y(n_688)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_682),
.Y(n_681)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_684),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_686),
.B(n_687),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_SL g690 ( 
.A(n_686),
.B(n_687),
.Y(n_690)
);

NOR3x1_ASAP7_75t_L g699 ( 
.A(n_700),
.B(n_702),
.C(n_703),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_706),
.Y(n_705)
);

INVx6_ASAP7_75t_L g706 ( 
.A(n_707),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_SL g708 ( 
.A1(n_709),
.A2(n_710),
.B(n_711),
.Y(n_708)
);


endmodule