module fake_jpeg_11955_n_187 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_2),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_19),
.B1(n_47),
.B2(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_58),
.B1(n_65),
.B2(n_67),
.Y(n_104)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_76),
.B1(n_62),
.B2(n_70),
.Y(n_100)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_95),
.C(n_97),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_74),
.B1(n_80),
.B2(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_64),
.B1(n_69),
.B2(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_79),
.Y(n_97)
);

OR2x6_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_73),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_60),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_78),
.B1(n_54),
.B2(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_105),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_83),
.B1(n_78),
.B2(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_112),
.B1(n_124),
.B2(n_126),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_72),
.B(n_63),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_122),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_98),
.B(n_95),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_27),
.B(n_45),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_105),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_24),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_8),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_56),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_7),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_146),
.B1(n_15),
.B2(n_33),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_8),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_9),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_147),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_36),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_26),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_11),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_13),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_34),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_154),
.C(n_165),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_129),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_35),
.B1(n_40),
.B2(n_44),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_162),
.Y(n_172)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_49),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_166),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_145),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_141),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_157),
.A3(n_158),
.B1(n_164),
.B2(n_151),
.C1(n_165),
.C2(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_173),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_178),
.B(n_179),
.C(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_175),
.B(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_160),
.C(n_170),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_180),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_179),
.C(n_168),
.Y(n_184)
);

AOI211xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_168),
.B(n_172),
.C(n_131),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_131),
.B(n_130),
.C(n_144),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_144),
.Y(n_187)
);


endmodule