module fake_jpeg_8214_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_20),
.B1(n_31),
.B2(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_41),
.B1(n_27),
.B2(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_34),
.B1(n_43),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_60),
.B1(n_25),
.B2(n_19),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_20),
.B1(n_31),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_62),
.B1(n_66),
.B2(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_57),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_31),
.B1(n_22),
.B2(n_24),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_68),
.Y(n_70)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_86),
.B1(n_49),
.B2(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_28),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_41),
.B1(n_25),
.B2(n_19),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_25),
.B1(n_19),
.B2(n_28),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_50),
.B1(n_32),
.B2(n_29),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_56),
.B1(n_53),
.B2(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_116),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_68),
.B1(n_63),
.B2(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_80),
.B1(n_79),
.B2(n_73),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_75),
.B(n_81),
.C(n_74),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_112),
.B(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_114),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_53),
.B(n_69),
.C(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_122),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_49),
.A3(n_63),
.B1(n_44),
.B2(n_57),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_71),
.B(n_74),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_67),
.B(n_50),
.C(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_45),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_119),
.B1(n_88),
.B2(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_0),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_23),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_148),
.C(n_122),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_126),
.B(n_141),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_0),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_136),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_89),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_112),
.B1(n_116),
.B2(n_57),
.Y(n_172)
);

OR2x2_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_147),
.B(n_111),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_98),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_159),
.C(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_107),
.B(n_113),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_157),
.B(n_167),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_117),
.B(n_115),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_124),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_99),
.C(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_134),
.B1(n_133),
.B2(n_114),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_141),
.B(n_127),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_136),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_127),
.C(n_134),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_174),
.B(n_131),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_173),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_112),
.B(n_116),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_180),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_189),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_158),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_193),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_191),
.B(n_192),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_141),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_132),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_132),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_171),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_167),
.B1(n_154),
.B2(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_197),
.B1(n_172),
.B2(n_129),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_140),
.B1(n_146),
.B2(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_171),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_203),
.B1(n_216),
.B2(n_176),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_153),
.B1(n_174),
.B2(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_218),
.B1(n_197),
.B2(n_196),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_157),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_183),
.C(n_193),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_160),
.B(n_162),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_215),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_160),
.C(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_172),
.B1(n_170),
.B2(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_199),
.B(n_105),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_236),
.B(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_183),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_237),
.C(n_242),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_184),
.C(n_194),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_202),
.A2(n_186),
.B1(n_182),
.B2(n_187),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_239),
.B1(n_205),
.B2(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_226),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_185),
.C(n_188),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_230),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_259),
.B1(n_254),
.B2(n_253),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_250),
.C(n_254),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_175),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_23),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_203),
.B1(n_180),
.B2(n_213),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_200),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_105),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_190),
.C(n_175),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_33),
.B(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_223),
.B(n_224),
.C(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_266),
.B1(n_268),
.B2(n_244),
.Y(n_275)
);

OAI311xp33_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_230),
.A3(n_172),
.B1(n_212),
.C1(n_135),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_247),
.B1(n_32),
.B2(n_10),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_273),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_249),
.B(n_255),
.C(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_271),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_172),
.B1(n_94),
.B2(n_87),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_8),
.C(n_15),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_94),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_247),
.B(n_87),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_280),
.B(n_281),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_266),
.B1(n_260),
.B2(n_11),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_285),
.B1(n_2),
.B2(n_4),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_87),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_7),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_9),
.B1(n_14),
.B2(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_1),
.C(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_264),
.C(n_3),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_7),
.B(n_13),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_12),
.B(n_14),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_9),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_288),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_280),
.B1(n_260),
.B2(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_277),
.C(n_274),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_6),
.B(n_13),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_6),
.Y(n_300)
);

AOI31xp67_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_260),
.A3(n_282),
.B(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_287),
.B(n_290),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_4),
.B(n_296),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_299),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_289),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_6),
.B(n_2),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_306),
.B(n_297),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_303),
.B(n_304),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_307),
.B(n_4),
.Y(n_311)
);


endmodule