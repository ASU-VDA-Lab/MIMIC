module real_aes_1267_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_838, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_837, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_838;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_837;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g185 ( .A(n_0), .B(n_159), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_1), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_2), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g150 ( .A(n_3), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_4), .B(n_143), .Y(n_212) );
NAND2xp33_ASAP7_75t_SL g255 ( .A(n_5), .B(n_149), .Y(n_255) );
INVx1_ASAP7_75t_L g247 ( .A(n_6), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_7), .B(n_217), .Y(n_505) );
INVx1_ASAP7_75t_L g486 ( .A(n_8), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_9), .Y(n_121) );
AND2x2_ASAP7_75t_L g210 ( .A(n_10), .B(n_167), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_11), .Y(n_569) );
INVx2_ASAP7_75t_L g165 ( .A(n_12), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
INVx1_ASAP7_75t_L g513 ( .A(n_14), .Y(n_513) );
AOI221x1_ASAP7_75t_L g250 ( .A1(n_15), .A2(n_152), .B1(n_251), .B2(n_253), .C(n_254), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_16), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g117 ( .A(n_17), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_18), .Y(n_802) );
INVx1_ASAP7_75t_L g511 ( .A(n_19), .Y(n_511) );
INVx1_ASAP7_75t_SL g523 ( .A(n_20), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_21), .B(n_144), .Y(n_501) );
AOI221xp5_ASAP7_75t_SL g174 ( .A1(n_22), .A2(n_43), .B1(n_143), .B2(n_152), .C(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_23), .A2(n_152), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_24), .B(n_159), .Y(n_215) );
AOI33xp33_ASAP7_75t_L g478 ( .A1(n_25), .A2(n_56), .A3(n_198), .B1(n_205), .B2(n_479), .B3(n_480), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_26), .A2(n_41), .B1(n_826), .B2(n_827), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_26), .Y(n_827) );
INVx1_ASAP7_75t_L g563 ( .A(n_27), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_28), .A2(n_125), .B1(n_126), .B2(n_132), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_28), .Y(n_132) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_29), .A2(n_93), .B(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g168 ( .A(n_29), .B(n_93), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_30), .B(n_161), .Y(n_160) );
INVxp67_ASAP7_75t_L g249 ( .A(n_31), .Y(n_249) );
AND2x2_ASAP7_75t_L g236 ( .A(n_32), .B(n_173), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_33), .B(n_196), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_34), .A2(n_152), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_35), .B(n_666), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g789 ( .A(n_35), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_36), .B(n_161), .Y(n_176) );
AND2x2_ASAP7_75t_L g149 ( .A(n_37), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g153 ( .A(n_37), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g204 ( .A(n_37), .Y(n_204) );
OR2x6_ASAP7_75t_L g115 ( .A(n_38), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_39), .A2(n_73), .B1(n_822), .B2(n_823), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_39), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_40), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_41), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_42), .B(n_196), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_44), .A2(n_127), .B1(n_128), .B2(n_129), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_44), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_45), .A2(n_181), .B1(n_217), .B2(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_46), .A2(n_85), .B1(n_152), .B2(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_47), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_48), .B(n_144), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_49), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_50), .B(n_159), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_51), .B(n_163), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_52), .B(n_144), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_53), .Y(n_498) );
AND2x2_ASAP7_75t_L g188 ( .A(n_54), .B(n_173), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_55), .B(n_173), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_57), .B(n_144), .Y(n_469) );
INVx1_ASAP7_75t_L g146 ( .A(n_58), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_58), .Y(n_156) );
AND2x2_ASAP7_75t_L g470 ( .A(n_59), .B(n_173), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_60), .A2(n_78), .B1(n_196), .B2(n_202), .C(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_61), .B(n_196), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_62), .B(n_143), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_63), .B(n_181), .Y(n_571) );
AOI21xp5_ASAP7_75t_SL g531 ( .A1(n_64), .A2(n_202), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g227 ( .A(n_65), .B(n_173), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_66), .B(n_161), .Y(n_186) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_67), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_68), .B(n_159), .Y(n_224) );
INVx1_ASAP7_75t_L g508 ( .A(n_69), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_70), .A2(n_152), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g467 ( .A(n_71), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_72), .B(n_161), .Y(n_216) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_73), .B(n_163), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_73), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_74), .A2(n_202), .B(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_75), .A2(n_97), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_75), .Y(n_130) );
INVx1_ASAP7_75t_L g148 ( .A(n_76), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_76), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_77), .B(n_196), .Y(n_481) );
AND2x2_ASAP7_75t_L g525 ( .A(n_79), .B(n_253), .Y(n_525) );
INVx1_ASAP7_75t_L g509 ( .A(n_80), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_81), .A2(n_202), .B(n_522), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_82), .A2(n_193), .B(n_202), .C(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_83), .A2(n_88), .B1(n_143), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_84), .B(n_143), .Y(n_225) );
INVx1_ASAP7_75t_L g118 ( .A(n_86), .Y(n_118) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_87), .B(n_253), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_89), .A2(n_202), .B1(n_476), .B2(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_90), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_91), .B(n_159), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_92), .A2(n_152), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g533 ( .A(n_94), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_95), .B(n_161), .Y(n_223) );
AND2x2_ASAP7_75t_L g482 ( .A(n_96), .B(n_253), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_97), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_98), .A2(n_561), .B(n_562), .C(n_564), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_99), .B(n_143), .Y(n_187) );
INVxp67_ASAP7_75t_L g252 ( .A(n_100), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_101), .B(n_161), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_102), .A2(n_152), .B(n_157), .Y(n_151) );
BUFx2_ASAP7_75t_L g812 ( .A(n_103), .Y(n_812) );
BUFx2_ASAP7_75t_SL g832 ( .A(n_103), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_104), .B(n_144), .Y(n_534) );
AOI21xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_122), .B(n_833), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g835 ( .A(n_109), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_119), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g806 ( .A(n_112), .Y(n_806) );
BUFx2_ASAP7_75t_R g817 ( .A(n_112), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_113), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_113), .B(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_SL g797 ( .A(n_113), .B(n_114), .Y(n_797) );
OR2x2_ASAP7_75t_L g810 ( .A(n_113), .B(n_115), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_115), .A2(n_124), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_813), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_133), .B(n_791), .C(n_793), .Y(n_123) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_124), .Y(n_799) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVxp33_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
OAI21xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_449), .B(n_451), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_SL g798 ( .A(n_135), .Y(n_798) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_341), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_269), .C(n_319), .Y(n_136) );
OAI211xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_189), .B(n_237), .C(n_258), .Y(n_137) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_169), .Y(n_138) );
AND2x2_ASAP7_75t_L g268 ( .A(n_139), .B(n_170), .Y(n_268) );
INVx1_ASAP7_75t_L g399 ( .A(n_139), .Y(n_399) );
NOR2x1p5_ASAP7_75t_L g431 ( .A(n_139), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g242 ( .A(n_140), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g290 ( .A(n_140), .Y(n_290) );
OR2x2_ASAP7_75t_L g294 ( .A(n_140), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_140), .B(n_172), .Y(n_306) );
OR2x2_ASAP7_75t_L g328 ( .A(n_140), .B(n_172), .Y(n_328) );
AND2x4_ASAP7_75t_L g334 ( .A(n_140), .B(n_298), .Y(n_334) );
OR2x2_ASAP7_75t_L g351 ( .A(n_140), .B(n_244), .Y(n_351) );
INVx1_ASAP7_75t_L g386 ( .A(n_140), .Y(n_386) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_140), .Y(n_408) );
OR2x2_ASAP7_75t_L g422 ( .A(n_140), .B(n_355), .Y(n_422) );
AND2x4_ASAP7_75t_SL g426 ( .A(n_140), .B(n_244), .Y(n_426) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_166), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_151), .B(n_163), .Y(n_141) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
AND2x6_ASAP7_75t_L g159 ( .A(n_145), .B(n_154), .Y(n_159) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g161 ( .A(n_147), .B(n_156), .Y(n_161) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_149), .Y(n_564) );
AND2x2_ASAP7_75t_L g155 ( .A(n_150), .B(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_150), .Y(n_199) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
BUFx3_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx2_ASAP7_75t_L g206 ( .A(n_154), .Y(n_206) );
AND2x4_ASAP7_75t_L g202 ( .A(n_155), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
INVxp67_ASAP7_75t_L g512 ( .A(n_159), .Y(n_512) );
INVxp67_ASAP7_75t_L g514 ( .A(n_161), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_162), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_162), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_162), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_162), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_162), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_162), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g476 ( .A(n_162), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_162), .A2(n_468), .B(n_486), .C(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_162), .A2(n_501), .B(n_502), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_162), .B(n_217), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_162), .A2(n_468), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_162), .A2(n_468), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_SL g193 ( .A(n_163), .Y(n_193) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_163), .A2(n_484), .B(n_488), .Y(n_483) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_165), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g217 ( .A(n_165), .B(n_168), .Y(n_217) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g378 ( .A(n_170), .B(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g425 ( .A(n_170), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_179), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
AND2x2_ASAP7_75t_L g288 ( .A(n_172), .B(n_179), .Y(n_288) );
INVx2_ASAP7_75t_L g295 ( .A(n_172), .Y(n_295) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_172), .Y(n_416) );
BUFx3_ASAP7_75t_L g432 ( .A(n_172), .Y(n_432) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_178), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_173), .Y(n_226) );
INVx2_ASAP7_75t_L g257 ( .A(n_179), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_179), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g355 ( .A(n_179), .B(n_295), .Y(n_355) );
INVx1_ASAP7_75t_L g373 ( .A(n_179), .Y(n_373) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_179), .Y(n_389) );
INVx1_ASAP7_75t_L g411 ( .A(n_179), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_179), .B(n_290), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_179), .B(n_244), .Y(n_448) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
INVx4_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_181), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_208), .Y(n_190) );
AND2x4_ASAP7_75t_L g262 ( .A(n_191), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_191), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_191), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g313 ( .A(n_191), .B(n_218), .Y(n_313) );
AND2x2_ASAP7_75t_L g323 ( .A(n_191), .B(n_219), .Y(n_323) );
OR2x2_ASAP7_75t_L g403 ( .A(n_191), .B(n_318), .Y(n_403) );
OAI322xp33_ASAP7_75t_L g433 ( .A1(n_191), .A2(n_346), .A3(n_385), .B1(n_418), .B2(n_434), .C1(n_435), .C2(n_436), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_191), .B(n_416), .Y(n_434) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
AOI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_207), .Y(n_192) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_193), .A2(n_474), .B(n_482), .Y(n_473) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_193), .A2(n_474), .B(n_482), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_201), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_196), .A2(n_202), .B1(n_246), .B2(n_248), .Y(n_245) );
INVx1_ASAP7_75t_L g572 ( .A(n_196), .Y(n_572) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_200), .Y(n_196) );
INVx1_ASAP7_75t_L g496 ( .A(n_197), .Y(n_496) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
OR2x6_ASAP7_75t_L g468 ( .A(n_198), .B(n_206), .Y(n_468) );
INVxp33_ASAP7_75t_L g479 ( .A(n_198), .Y(n_479) );
INVx1_ASAP7_75t_L g497 ( .A(n_200), .Y(n_497) );
INVxp67_ASAP7_75t_L g570 ( .A(n_202), .Y(n_570) );
NOR2x1p5_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g480 ( .A(n_205), .Y(n_480) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_208), .A2(n_380), .B1(n_384), .B2(n_387), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_208), .A2(n_440), .B(n_441), .C(n_444), .Y(n_439) );
AND2x4_ASAP7_75t_SL g208 ( .A(n_209), .B(n_218), .Y(n_208) );
AND2x4_ASAP7_75t_L g261 ( .A(n_209), .B(n_229), .Y(n_261) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
INVx5_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
INVx2_ASAP7_75t_L g286 ( .A(n_209), .Y(n_286) );
AND2x2_ASAP7_75t_L g309 ( .A(n_209), .B(n_219), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_209), .B(n_228), .Y(n_338) );
OR2x2_ASAP7_75t_L g347 ( .A(n_209), .B(n_267), .Y(n_347) );
OR2x2_ASAP7_75t_L g362 ( .A(n_209), .B(n_276), .Y(n_362) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_217), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_217), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_217), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_217), .B(n_252), .Y(n_251) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_217), .B(n_255), .C(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_217), .A2(n_531), .B(n_535), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_218), .B(n_238), .Y(n_237) );
INVx3_ASAP7_75t_SL g346 ( .A(n_218), .Y(n_346) );
AND2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_277), .Y(n_369) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
AND2x2_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g280 ( .A(n_219), .B(n_229), .Y(n_280) );
INVx1_ASAP7_75t_L g284 ( .A(n_219), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_219), .B(n_229), .Y(n_318) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_219), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_219), .B(n_277), .Y(n_393) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_227), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_226), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_226), .A2(n_230), .B(n_236), .Y(n_276) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_226), .A2(n_519), .B(n_525), .Y(n_518) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
AND2x2_ASAP7_75t_L g383 ( .A(n_229), .B(n_267), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x6_ASAP7_75t_SL g447 ( .A(n_240), .B(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_241), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_241), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g395 ( .A(n_241), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_242), .A2(n_304), .B1(n_307), .B2(n_314), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_243), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_243), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_243), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_243), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_257), .Y(n_243) );
AND2x2_ASAP7_75t_L g289 ( .A(n_244), .B(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_244), .A2(n_305), .B1(n_357), .B2(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g364 ( .A(n_244), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_244), .B(n_358), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_244), .B(n_288), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_244), .B(n_295), .Y(n_437) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
INVx3_ASAP7_75t_L g462 ( .A(n_253), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_253), .A2(n_462), .B1(n_560), .B2(n_565), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_256), .A2(n_468), .B1(n_508), .B2(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_256), .B(n_563), .Y(n_562) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B(n_268), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
NAND4xp25_ASAP7_75t_SL g307 ( .A(n_260), .B(n_308), .C(n_310), .D(n_312), .Y(n_307) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_261), .B(n_368), .Y(n_397) );
AND2x2_ASAP7_75t_L g424 ( .A(n_261), .B(n_262), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_261), .B(n_284), .Y(n_435) );
INVx1_ASAP7_75t_L g300 ( .A(n_262), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_262), .A2(n_325), .B1(n_336), .B2(n_339), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_262), .B(n_275), .C(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_262), .B(n_277), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_262), .B(n_285), .Y(n_428) );
AND2x2_ASAP7_75t_L g360 ( .A(n_263), .B(n_267), .Y(n_360) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_263), .Y(n_421) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g316 ( .A(n_265), .Y(n_316) );
INVx1_ASAP7_75t_L g406 ( .A(n_266), .Y(n_406) );
AND2x2_ASAP7_75t_L g413 ( .A(n_266), .B(n_277), .Y(n_413) );
BUFx2_ASAP7_75t_L g368 ( .A(n_267), .Y(n_368) );
NAND3xp33_ASAP7_75t_SL g269 ( .A(n_270), .B(n_291), .C(n_303), .Y(n_269) );
OAI31xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_278), .A3(n_281), .B(n_287), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_325), .B1(n_329), .B2(n_330), .Y(n_324) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g310 ( .A(n_273), .B(n_311), .Y(n_310) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_273), .B(n_337), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_274), .A2(n_376), .B(n_406), .C(n_407), .Y(n_405) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_275), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_276), .B(n_284), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_309), .Y(n_329) );
AND2x2_ASAP7_75t_L g446 ( .A(n_279), .B(n_368), .Y(n_446) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g302 ( .A(n_280), .B(n_286), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_360), .Y(n_377) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_286), .B(n_360), .Y(n_366) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g358 ( .A(n_288), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_289), .B(n_389), .Y(n_388) );
AOI32xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_299), .A3(n_300), .B1(n_301), .B2(n_837), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_292), .A2(n_377), .B1(n_413), .B2(n_414), .C(n_417), .Y(n_412) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g305 ( .A(n_297), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g410 ( .A(n_298), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_299), .B(n_321), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_301), .A2(n_344), .B1(n_348), .B2(n_352), .C(n_356), .Y(n_343) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_306), .A2(n_320), .B(n_324), .C(n_335), .Y(n_319) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g417 ( .A1(n_312), .A2(n_322), .A3(n_371), .B1(n_418), .B2(n_419), .C1(n_420), .C2(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_315), .A2(n_445), .B(n_447), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_321), .A2(n_402), .B(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g443 ( .A(n_328), .B(n_409), .Y(n_443) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_334), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g418 ( .A(n_334), .Y(n_418) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_375), .A3(n_377), .B(n_378), .Y(n_374) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_400), .Y(n_341) );
NAND5xp2_ASAP7_75t_L g342 ( .A(n_343), .B(n_363), .C(n_374), .D(n_379), .E(n_390), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_346), .A2(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g414 ( .A(n_350), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_367), .C(n_370), .Y(n_363) );
INVxp33_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g392 ( .A(n_368), .B(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_371), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g442 ( .A(n_383), .Y(n_442) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_392), .A2(n_397), .B(n_398), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .C(n_423), .D(n_439), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_410), .B(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_433), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g792 ( .A(n_451), .Y(n_792) );
INVx2_ASAP7_75t_L g819 ( .A(n_452), .Y(n_819) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_786), .Y(n_452) );
NOR4xp25_ASAP7_75t_L g453 ( .A(n_454), .B(n_665), .C(n_689), .D(n_755), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_454), .A2(n_689), .B1(n_789), .B2(n_838), .Y(n_790) );
NAND3x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_617), .C(n_651), .Y(n_454) );
NOR3x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_576), .C(n_596), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_551), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_489), .B1(n_540), .B2(n_548), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_471), .Y(n_458) );
AND2x2_ASAP7_75t_L g715 ( .A(n_459), .B(n_645), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_459), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_459), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_459), .B(n_585), .Y(n_774) );
OR2x2_ASAP7_75t_L g784 ( .A(n_459), .B(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g605 ( .A(n_460), .B(n_542), .Y(n_605) );
AND2x4_ASAP7_75t_L g633 ( .A(n_460), .B(n_547), .Y(n_633) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g581 ( .A(n_461), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_461), .B(n_473), .Y(n_671) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_461), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_461), .B(n_558), .Y(n_708) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_470), .Y(n_461) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_462), .A2(n_463), .B(n_470), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g503 ( .A(n_468), .Y(n_503) );
INVxp67_ASAP7_75t_L g561 ( .A(n_468), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_471), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g779 ( .A(n_471), .B(n_616), .Y(n_779) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g769 ( .A(n_472), .B(n_708), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
INVx2_ASAP7_75t_L g547 ( .A(n_473), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_475), .B(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
INVx2_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_483), .Y(n_582) );
INVx1_ASAP7_75t_L g595 ( .A(n_483), .Y(n_595) );
INVxp67_ASAP7_75t_L g614 ( .A(n_483), .Y(n_614) );
AND2x4_ASAP7_75t_L g645 ( .A(n_483), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_526), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_516), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g687 ( .A(n_492), .B(n_674), .Y(n_687) );
AND2x2_ASAP7_75t_L g711 ( .A(n_492), .B(n_527), .Y(n_711) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
INVx2_ASAP7_75t_L g539 ( .A(n_493), .Y(n_539) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
INVx1_ASAP7_75t_L g611 ( .A(n_493), .Y(n_611) );
AND2x4_ASAP7_75t_L g620 ( .A(n_493), .B(n_538), .Y(n_620) );
AND2x2_ASAP7_75t_L g676 ( .A(n_493), .B(n_528), .Y(n_676) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_499), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .C(n_498), .Y(n_495) );
INVx3_ASAP7_75t_L g538 ( .A(n_504), .Y(n_538) );
AND2x2_ASAP7_75t_L g550 ( .A(n_504), .B(n_518), .Y(n_550) );
INVx2_ASAP7_75t_L g589 ( .A(n_504), .Y(n_589) );
NOR2x1_ASAP7_75t_SL g602 ( .A(n_504), .B(n_528), .Y(n_602) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .B(n_515), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g704 ( .A(n_516), .Y(n_704) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g627 ( .A(n_517), .Y(n_627) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_518), .Y(n_601) );
AND2x2_ASAP7_75t_L g609 ( .A(n_518), .B(n_538), .Y(n_609) );
INVx1_ASAP7_75t_L g649 ( .A(n_518), .Y(n_649) );
INVx1_ASAP7_75t_L g674 ( .A(n_518), .Y(n_674) );
OR2x2_ASAP7_75t_L g735 ( .A(n_518), .B(n_528), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
OA211x2_ASAP7_75t_L g756 ( .A1(n_526), .A2(n_757), .B(n_759), .C(n_766), .Y(n_756) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
AND2x2_ASAP7_75t_L g677 ( .A(n_527), .B(n_550), .Y(n_677) );
AND2x2_ASAP7_75t_SL g695 ( .A(n_527), .B(n_537), .Y(n_695) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
INVx2_ASAP7_75t_L g591 ( .A(n_528), .Y(n_591) );
AND2x4_ASAP7_75t_L g654 ( .A(n_528), .B(n_611), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_528), .B(n_650), .Y(n_705) );
AND2x2_ASAP7_75t_L g748 ( .A(n_528), .B(n_589), .Y(n_748) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_537), .B(n_649), .Y(n_742) );
AND2x2_ASAP7_75t_L g762 ( .A(n_537), .B(n_585), .Y(n_762) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g650 ( .A(n_538), .Y(n_650) );
INVx1_ASAP7_75t_L g624 ( .A(n_539), .Y(n_624) );
NOR2xp67_ASAP7_75t_SL g540 ( .A(n_541), .B(n_544), .Y(n_540) );
INVx1_ASAP7_75t_L g718 ( .A(n_541), .Y(n_718) );
NOR2xp67_ASAP7_75t_L g765 ( .A(n_541), .B(n_719), .Y(n_765) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g738 ( .A(n_543), .B(n_580), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_544), .A2(n_727), .B(n_730), .C(n_739), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_544), .A2(n_764), .B(n_771), .C(n_775), .Y(n_770) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g655 ( .A(n_545), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g574 ( .A(n_546), .Y(n_574) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_546), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g630 ( .A(n_546), .B(n_580), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g740 ( .A(n_546), .B(n_580), .Y(n_740) );
AND2x2_ASAP7_75t_L g613 ( .A(n_547), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g664 ( .A(n_547), .Y(n_664) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x4_ASAP7_75t_SL g553 ( .A(n_549), .B(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g610 ( .A(n_549), .B(n_611), .Y(n_610) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_549), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g658 ( .A(n_549), .B(n_659), .Y(n_658) );
NOR2xp67_ASAP7_75t_SL g741 ( .A(n_549), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_550), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_SL g781 ( .A(n_550), .B(n_623), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx2_ASAP7_75t_SL g749 ( .A(n_555), .Y(n_749) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_573), .Y(n_555) );
INVx3_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
AND2x2_ASAP7_75t_L g693 ( .A(n_556), .B(n_684), .Y(n_693) );
AND2x2_ASAP7_75t_L g751 ( .A(n_556), .B(n_633), .Y(n_751) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g580 ( .A(n_558), .Y(n_580) );
INVx1_ASAP7_75t_L g616 ( .A(n_558), .Y(n_616) );
INVx1_ASAP7_75t_L g636 ( .A(n_558), .Y(n_636) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_566), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_566) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVxp67_ASAP7_75t_L g719 ( .A(n_573), .Y(n_719) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_575), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g646 ( .A(n_575), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_583), .B1(n_586), .B2(n_592), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g593 ( .A(n_579), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g604 ( .A(n_579), .Y(n_604) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g653 ( .A(n_584), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g673 ( .A(n_588), .B(n_674), .Y(n_673) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g681 ( .A(n_589), .Y(n_681) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g729 ( .A(n_591), .B(n_620), .Y(n_729) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_593), .A2(n_687), .B(n_688), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_603), .B(n_606), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g652 ( .A(n_602), .B(n_626), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_603), .A2(n_710), .B1(n_712), .B2(n_714), .Y(n_709) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_612), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_SL g659 ( .A(n_609), .Y(n_659) );
AND2x2_ASAP7_75t_L g688 ( .A(n_610), .B(n_626), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_610), .B(n_648), .Y(n_720) );
AND2x2_ASAP7_75t_L g724 ( .A(n_610), .B(n_681), .Y(n_724) );
OAI21xp5_ASAP7_75t_SL g668 ( .A1(n_612), .A2(n_669), .B(n_673), .Y(n_668) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g629 ( .A(n_613), .B(n_630), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_613), .B(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g698 ( .A(n_616), .Y(n_698) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_641), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_628), .B1(n_631), .B2(n_637), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx4_ASAP7_75t_L g640 ( .A(n_620), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_620), .B(n_626), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_620), .B(n_773), .Y(n_772) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_623), .A2(n_647), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g746 ( .A(n_623), .B(n_648), .Y(n_746) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g728 ( .A(n_625), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g764 ( .A(n_626), .B(n_748), .Y(n_764) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g644 ( .A(n_630), .B(n_645), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_630), .B(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_SL g641 ( .A1(n_631), .A2(n_642), .B1(n_643), .B2(n_647), .Y(n_641) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g758 ( .A(n_635), .B(n_645), .Y(n_758) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g656 ( .A(n_636), .Y(n_656) );
AND2x2_ASAP7_75t_L g682 ( .A(n_636), .B(n_645), .Y(n_682) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_638), .B(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_639), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g733 ( .A(n_640), .Y(n_733) );
INVx1_ASAP7_75t_L g745 ( .A(n_642), .Y(n_745) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_644), .A2(n_688), .B1(n_767), .B2(n_768), .Y(n_766) );
AND2x2_ASAP7_75t_L g683 ( .A(n_645), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g754 ( .A(n_645), .B(n_707), .Y(n_754) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI211xp5_ASAP7_75t_SL g657 ( .A1(n_648), .A2(n_658), .B(n_660), .C(n_661), .Y(n_657) );
AND2x2_ASAP7_75t_SL g767 ( .A(n_648), .B(n_654), .Y(n_767) );
AND2x4_ASAP7_75t_SL g648 ( .A(n_649), .B(n_650), .Y(n_648) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_649), .Y(n_701) );
O2A1O1Ixp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_655), .C(n_657), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_652), .A2(n_680), .B1(n_682), .B2(n_683), .Y(n_679) );
INVx2_ASAP7_75t_L g660 ( .A(n_654), .Y(n_660) );
AND2x2_ASAP7_75t_L g680 ( .A(n_654), .B(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_654), .Y(n_747) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g788 ( .A(n_666), .Y(n_788) );
NOR2x1_ASAP7_75t_SL g666 ( .A(n_667), .B(n_678), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_675), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_669), .A2(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g699 ( .A(n_671), .Y(n_699) );
INVx1_ASAP7_75t_L g775 ( .A(n_672), .Y(n_775) );
AND2x2_ASAP7_75t_L g713 ( .A(n_676), .B(n_701), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_677), .B(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_686), .Y(n_678) );
AND2x2_ASAP7_75t_L g780 ( .A(n_682), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_725), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_709), .C(n_716), .Y(n_690) );
OAI222xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B1(n_696), .B2(n_700), .C1(n_702), .C2(n_706), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g752 ( .A(n_711), .Y(n_752) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NOR2xp67_ASAP7_75t_SL g725 ( .A(n_726), .B(n_743), .Y(n_725) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_733), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g785 ( .A(n_738), .Y(n_785) );
NAND2xp33_ASAP7_75t_SL g739 ( .A(n_740), .B(n_741), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_749), .B1(n_750), .B2(n_752), .C(n_753), .Y(n_743) );
NOR4xp25_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .C(n_747), .D(n_748), .Y(n_744) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_755), .A2(n_788), .B(n_789), .Y(n_787) );
NAND4xp75_ASAP7_75t_L g755 ( .A(n_756), .B(n_770), .C(n_776), .D(n_782), .Y(n_755) );
INVx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_760), .B(n_765), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_790), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_799), .B(n_800), .Y(n_793) );
INVxp33_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2x1_ASAP7_75t_SL g795 ( .A(n_796), .B(n_798), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
OR3x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_807), .C(n_811), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_801), .A2(n_815), .B(n_818), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_829), .Y(n_813) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_824), .B1(n_825), .B2(n_828), .Y(n_820) );
INVx1_ASAP7_75t_L g828 ( .A(n_821), .Y(n_828) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
CKINVDCx11_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
endmodule