module real_aes_7438_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_698, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_698;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_668;
wire n_237;
A2O1A1Ixp33_ASAP7_75t_SL g152 ( .A1(n_0), .A2(n_153), .B(n_154), .C(n_158), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_1), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_2), .B(n_147), .Y(n_160) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_4), .B(n_132), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g428 ( .A1(n_5), .A2(n_121), .B(n_138), .C(n_429), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_6), .A2(n_141), .B(n_450), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_7), .A2(n_141), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_8), .B(n_147), .Y(n_456) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_9), .A2(n_113), .B(n_200), .Y(n_199) );
AND2x6_ASAP7_75t_L g138 ( .A(n_10), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_11), .A2(n_121), .B(n_138), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g421 ( .A(n_12), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_13), .B(n_40), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_14), .B(n_157), .Y(n_431) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_16), .B(n_132), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_17), .A2(n_133), .B(n_440), .C(n_442), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_18), .B(n_147), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_19), .A2(n_99), .B1(n_670), .B2(n_679), .C1(n_688), .C2(n_694), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g681 ( .A1(n_19), .A2(n_662), .B1(n_682), .B2(n_683), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_19), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_20), .B(n_190), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_21), .A2(n_121), .B(n_184), .C(n_189), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_22), .A2(n_156), .B(n_208), .C(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_23), .B(n_157), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_24), .B(n_157), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_25), .Y(n_459) );
INVx1_ASAP7_75t_L g471 ( .A(n_26), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_27), .A2(n_121), .B(n_189), .C(n_203), .Y(n_202) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_28), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_29), .Y(n_427) );
INVx1_ASAP7_75t_L g488 ( .A(n_30), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_31), .A2(n_141), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g123 ( .A(n_32), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_33), .A2(n_136), .B(n_168), .C(n_169), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_34), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_35), .A2(n_156), .B(n_453), .C(n_455), .Y(n_452) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_37), .B(n_205), .Y(n_204) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_38), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_39), .A2(n_121), .B(n_189), .C(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_41), .A2(n_158), .B(n_419), .C(n_420), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_42), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_43), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_44), .B(n_132), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_45), .B(n_141), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_46), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_48), .A2(n_136), .B(n_168), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_49), .Y(n_685) );
INVx1_ASAP7_75t_L g155 ( .A(n_50), .Y(n_155) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_100), .B1(n_661), .B2(n_665), .C1(n_666), .C2(n_669), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_51), .Y(n_665) );
INVx1_ASAP7_75t_L g230 ( .A(n_52), .Y(n_230) );
INVx1_ASAP7_75t_L g409 ( .A(n_53), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_54), .B(n_141), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
CKINVDCx14_ASAP7_75t_R g417 ( .A(n_56), .Y(n_417) );
INVx1_ASAP7_75t_L g139 ( .A(n_57), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_58), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_59), .B(n_147), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_60), .A2(n_128), .B(n_188), .C(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g117 ( .A(n_61), .Y(n_117) );
INVx1_ASAP7_75t_SL g454 ( .A(n_62), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_63), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_64), .B(n_132), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_65), .B(n_147), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_66), .B(n_133), .Y(n_219) );
INVx1_ASAP7_75t_L g462 ( .A(n_67), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_68), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_69), .B(n_172), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g120 ( .A1(n_70), .A2(n_121), .B(n_126), .C(n_136), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_71), .Y(n_244) );
INVx1_ASAP7_75t_L g674 ( .A(n_72), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_73), .A2(n_141), .B(n_416), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_74), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_75), .A2(n_141), .B(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_76), .A2(n_182), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g438 ( .A(n_77), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_78), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_79), .B(n_171), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_80), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_81), .A2(n_141), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g441 ( .A(n_82), .Y(n_441) );
INVx2_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
INVx1_ASAP7_75t_L g430 ( .A(n_84), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_85), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_86), .B(n_157), .Y(n_220) );
OR2x2_ASAP7_75t_L g102 ( .A(n_87), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g399 ( .A(n_87), .Y(n_399) );
OR2x2_ASAP7_75t_L g678 ( .A(n_87), .B(n_668), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_88), .A2(n_121), .B(n_136), .C(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_89), .B(n_141), .Y(n_166) );
INVx1_ASAP7_75t_L g170 ( .A(n_90), .Y(n_170) );
INVxp67_ASAP7_75t_L g247 ( .A(n_91), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_92), .B(n_113), .Y(n_422) );
INVx1_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
INVx1_ASAP7_75t_L g215 ( .A(n_94), .Y(n_215) );
INVx2_ASAP7_75t_L g412 ( .A(n_95), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_96), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g232 ( .A(n_97), .B(n_175), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_106), .B1(n_397), .B2(n_400), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_101), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x2_ASAP7_75t_L g398 ( .A(n_103), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g668 ( .A(n_103), .Y(n_668) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx2_ASAP7_75t_L g662 ( .A(n_106), .Y(n_662) );
NAND2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_340), .Y(n_106) );
AND4x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_280), .C(n_295), .D(n_320), .Y(n_107) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_253), .Y(n_108) );
OAI21xp33_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_161), .B(n_233), .Y(n_109) );
AND2x2_ASAP7_75t_L g283 ( .A(n_110), .B(n_179), .Y(n_283) );
AND2x2_ASAP7_75t_L g296 ( .A(n_110), .B(n_178), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_110), .B(n_162), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_110), .Y(n_350) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_146), .Y(n_110) );
INVx2_ASAP7_75t_L g267 ( .A(n_111), .Y(n_267) );
BUFx2_ASAP7_75t_L g294 ( .A(n_111), .Y(n_294) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_144), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_112), .B(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_112), .B(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_112), .A2(n_214), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_112), .B(n_434), .Y(n_433) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_112), .A2(n_458), .B(n_464), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_112), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_113), .A2(n_201), .B(n_202), .Y(n_200) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_113), .Y(n_241) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g223 ( .A(n_114), .Y(n_223) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_115), .B(n_116), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_140), .Y(n_119) );
INVx5_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
AND2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
BUFx3_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
INVx1_ASAP7_75t_L g209 ( .A(n_123), .Y(n_209) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_125), .Y(n_130) );
INVx3_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
AND2x2_ASAP7_75t_L g142 ( .A(n_125), .B(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx1_ASAP7_75t_L g205 ( .A(n_125), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_131), .C(n_134), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_129), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_129), .B(n_441), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_129), .A2(n_132), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
INVx2_ASAP7_75t_L g153 ( .A(n_132), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_132), .B(n_247), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_132), .A2(n_187), .B(n_471), .C(n_472), .Y(n_470) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_133), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g455 ( .A(n_135), .Y(n_455) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_SL g149 ( .A1(n_137), .A2(n_150), .B(n_151), .C(n_152), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_137), .A2(n_151), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g408 ( .A1(n_137), .A2(n_151), .B(n_409), .C(n_410), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_SL g416 ( .A1(n_137), .A2(n_151), .B(n_417), .C(n_418), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g437 ( .A1(n_137), .A2(n_151), .B(n_438), .C(n_439), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_137), .A2(n_151), .B(n_451), .C(n_452), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_137), .A2(n_151), .B(n_485), .C(n_486), .Y(n_484) );
INVx4_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g141 ( .A(n_138), .B(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_138), .B(n_142), .Y(n_216) );
BUFx2_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx1_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
AND2x2_ASAP7_75t_L g234 ( .A(n_146), .B(n_179), .Y(n_234) );
INVx2_ASAP7_75t_L g250 ( .A(n_146), .Y(n_250) );
AND2x2_ASAP7_75t_L g259 ( .A(n_146), .B(n_178), .Y(n_259) );
AND2x2_ASAP7_75t_L g338 ( .A(n_146), .B(n_267), .Y(n_338) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_160), .Y(n_146) );
INVx2_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_156), .B(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g419 ( .A(n_157), .Y(n_419) );
INVx2_ASAP7_75t_L g432 ( .A(n_158), .Y(n_432) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
INVx1_ASAP7_75t_L g442 ( .A(n_159), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_195), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_162), .B(n_265), .Y(n_303) );
INVx1_ASAP7_75t_L g391 ( .A(n_162), .Y(n_391) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_178), .Y(n_162) );
AND2x2_ASAP7_75t_L g249 ( .A(n_163), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g263 ( .A(n_163), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_163), .Y(n_292) );
OR2x2_ASAP7_75t_L g324 ( .A(n_163), .B(n_266), .Y(n_324) );
AND2x2_ASAP7_75t_L g332 ( .A(n_163), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g365 ( .A(n_163), .B(n_334), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_163), .B(n_234), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_163), .B(n_294), .Y(n_390) );
AND2x2_ASAP7_75t_L g396 ( .A(n_163), .B(n_283), .Y(n_396) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx2_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
AND2x2_ASAP7_75t_L g286 ( .A(n_164), .B(n_266), .Y(n_286) );
AND2x2_ASAP7_75t_L g319 ( .A(n_164), .B(n_279), .Y(n_319) );
AND2x2_ASAP7_75t_L g339 ( .A(n_164), .B(n_179), .Y(n_339) );
AND2x2_ASAP7_75t_L g373 ( .A(n_164), .B(n_239), .Y(n_373) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_176), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_175), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_173), .C(n_174), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_171), .A2(n_174), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp5_ASAP7_75t_L g429 ( .A1(n_171), .A2(n_430), .B(n_431), .C(n_432), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_171), .A2(n_432), .B(n_462), .C(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_175), .A2(n_227), .B(n_228), .Y(n_226) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_175), .A2(n_415), .B(n_422), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_175), .A2(n_216), .B(n_468), .C(n_469), .Y(n_467) );
AND2x4_ASAP7_75t_L g279 ( .A(n_178), .B(n_250), .Y(n_279) );
AND2x2_ASAP7_75t_L g290 ( .A(n_178), .B(n_286), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_178), .B(n_266), .Y(n_329) );
INVx2_ASAP7_75t_L g344 ( .A(n_178), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_178), .B(n_278), .Y(n_367) );
AND2x2_ASAP7_75t_L g386 ( .A(n_178), .B(n_338), .Y(n_386) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_179), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_179), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g334 ( .A(n_179), .B(n_250), .Y(n_334) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_192), .Y(n_179) );
AOI21xp5_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_183), .B(n_190), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_188), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_191), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AO21x2_ASAP7_75t_L g425 ( .A1(n_194), .A2(n_426), .B(n_433), .Y(n_425) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_210), .Y(n_196) );
AND2x2_ASAP7_75t_L g257 ( .A(n_197), .B(n_240), .Y(n_257) );
INVx1_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_198), .B(n_213), .Y(n_237) );
OR2x2_ASAP7_75t_L g270 ( .A(n_198), .B(n_240), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_198), .B(n_240), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_198), .B(n_239), .Y(n_302) );
AND2x2_ASAP7_75t_L g354 ( .A(n_198), .B(n_212), .Y(n_354) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_199), .B(n_224), .Y(n_262) );
AND2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_213), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B(n_207), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_207), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_210), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g288 ( .A(n_211), .B(n_270), .Y(n_288) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_224), .Y(n_211) );
OAI322xp33_ASAP7_75t_L g253 ( .A1(n_212), .A2(n_254), .A3(n_258), .B1(n_260), .B2(n_263), .C1(n_268), .C2(n_276), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_212), .B(n_239), .Y(n_261) );
OR2x2_ASAP7_75t_L g271 ( .A(n_212), .B(n_225), .Y(n_271) );
AND2x2_ASAP7_75t_L g273 ( .A(n_212), .B(n_225), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_212), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_212), .B(n_240), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_212), .B(n_369), .Y(n_368) );
INVx5_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_213), .B(n_257), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_216), .A2(n_427), .B(n_428), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_216), .A2(n_459), .B(n_460), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g482 ( .A(n_223), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_224), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g251 ( .A(n_224), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_224), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g313 ( .A(n_224), .B(n_240), .Y(n_313) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_224), .A2(n_342), .B(n_345), .C(n_357), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_224), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g379 ( .A(n_224), .B(n_354), .Y(n_379) );
INVx5_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g307 ( .A(n_225), .B(n_240), .Y(n_307) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_225), .Y(n_316) );
AND2x2_ASAP7_75t_L g356 ( .A(n_225), .B(n_354), .Y(n_356) );
AND2x2_ASAP7_75t_SL g387 ( .A(n_225), .B(n_257), .Y(n_387) );
AND2x2_ASAP7_75t_L g394 ( .A(n_225), .B(n_353), .Y(n_394) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_249), .B2(n_251), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_234), .B(n_256), .Y(n_304) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g252 ( .A(n_237), .Y(n_252) );
OR2x2_ASAP7_75t_L g312 ( .A(n_237), .B(n_313), .Y(n_312) );
OAI221xp5_ASAP7_75t_SL g360 ( .A1(n_237), .A2(n_361), .B1(n_363), .B2(n_364), .C(n_366), .Y(n_360) );
INVx2_ASAP7_75t_L g299 ( .A(n_238), .Y(n_299) );
AND2x2_ASAP7_75t_L g272 ( .A(n_239), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g362 ( .A(n_239), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_239), .B(n_354), .Y(n_375) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVxp67_ASAP7_75t_L g317 ( .A(n_240), .Y(n_317) );
AND2x2_ASAP7_75t_L g353 ( .A(n_240), .B(n_354), .Y(n_353) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_248), .Y(n_240) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_241), .A2(n_407), .B(n_413), .Y(n_406) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_241), .A2(n_436), .B(n_443), .Y(n_435) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_241), .A2(n_449), .B(n_456), .Y(n_448) );
AND2x2_ASAP7_75t_L g355 ( .A(n_249), .B(n_294), .Y(n_355) );
AND2x2_ASAP7_75t_L g265 ( .A(n_250), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_250), .B(n_323), .Y(n_322) );
NOR2xp33_ASAP7_75t_SL g336 ( .A(n_252), .B(n_299), .Y(n_336) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g342 ( .A(n_255), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OR2x2_ASAP7_75t_L g328 ( .A(n_256), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g393 ( .A(n_256), .B(n_338), .Y(n_393) );
INVx2_ASAP7_75t_L g326 ( .A(n_257), .Y(n_326) );
NAND4xp25_ASAP7_75t_SL g389 ( .A(n_258), .B(n_390), .C(n_391), .D(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_259), .B(n_323), .Y(n_358) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_SL g395 ( .A(n_262), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_SL g357 ( .A1(n_263), .A2(n_326), .B(n_330), .C(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g352 ( .A(n_265), .B(n_344), .Y(n_352) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_266), .Y(n_278) );
INVx1_ASAP7_75t_L g333 ( .A(n_266), .Y(n_333) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
AOI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B(n_272), .C(n_274), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_269), .B(n_273), .Y(n_289) );
OAI322xp33_ASAP7_75t_SL g327 ( .A1(n_269), .A2(n_328), .A3(n_330), .B1(n_331), .B2(n_335), .C1(n_336), .C2(n_337), .Y(n_327) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g349 ( .A(n_271), .B(n_275), .Y(n_349) );
INVx1_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
INVx1_ASAP7_75t_SL g348 ( .A(n_275), .Y(n_348) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_287), .B1(n_289), .B2(n_290), .C1(n_291), .C2(n_698), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_284), .Y(n_281) );
OAI322xp33_ASAP7_75t_L g370 ( .A1(n_282), .A2(n_344), .A3(n_349), .B1(n_371), .B2(n_372), .C1(n_374), .C2(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_283), .A2(n_297), .B1(n_321), .B2(n_325), .C(n_327), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OAI222xp33_ASAP7_75t_L g300 ( .A1(n_288), .A2(n_301), .B1(n_303), .B2(n_304), .C1(n_305), .C2(n_308), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_290), .A2(n_297), .B1(n_367), .B2(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_300), .C(n_311), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_297), .A2(n_334), .B(n_377), .C(n_380), .Y(n_376) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g369 ( .A(n_302), .Y(n_369) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_309), .B(n_334), .Y(n_363) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B(n_318), .Y(n_311) );
OAI221xp5_ASAP7_75t_SL g380 ( .A1(n_312), .A2(n_381), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_380) );
INVxp33_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_316), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_323), .B(n_334), .Y(n_374) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g385 ( .A(n_338), .B(n_344), .Y(n_385) );
AND4x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_359), .C(n_376), .D(n_388), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_351), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_355), .B2(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
INVx1_ASAP7_75t_SL g371 ( .A(n_356), .Y(n_371) );
NOR2xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_370), .Y(n_359) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_372), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_379), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx6_ASAP7_75t_L g663 ( .A(n_398), .Y(n_663) );
NOR2x2_ASAP7_75t_L g667 ( .A(n_399), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g664 ( .A(n_401), .Y(n_664) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_587), .Y(n_401) );
NOR4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_529), .C(n_559), .D(n_569), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_444), .B(n_492), .C(n_519), .Y(n_403) );
OAI222xp33_ASAP7_75t_L g614 ( .A1(n_404), .A2(n_534), .B1(n_615), .B2(n_616), .C1(n_617), .C2(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_423), .Y(n_404) );
AOI33xp33_ASAP7_75t_L g540 ( .A1(n_405), .A2(n_527), .A3(n_528), .B1(n_541), .B2(n_546), .B3(n_548), .Y(n_540) );
OAI211xp5_ASAP7_75t_SL g597 ( .A1(n_405), .A2(n_598), .B(n_600), .C(n_602), .Y(n_597) );
OR2x2_ASAP7_75t_L g613 ( .A(n_405), .B(n_599), .Y(n_613) );
INVx1_ASAP7_75t_L g646 ( .A(n_405), .Y(n_646) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_414), .Y(n_405) );
INVx2_ASAP7_75t_L g523 ( .A(n_406), .Y(n_523) );
AND2x2_ASAP7_75t_L g539 ( .A(n_406), .B(n_435), .Y(n_539) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_406), .Y(n_574) );
AND2x2_ASAP7_75t_L g603 ( .A(n_406), .B(n_414), .Y(n_603) );
INVx2_ASAP7_75t_L g503 ( .A(n_414), .Y(n_503) );
BUFx3_ASAP7_75t_L g511 ( .A(n_414), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_414), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g522 ( .A(n_414), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_414), .B(n_424), .Y(n_551) );
AND2x2_ASAP7_75t_L g620 ( .A(n_414), .B(n_554), .Y(n_620) );
INVx2_ASAP7_75t_SL g514 ( .A(n_423), .Y(n_514) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_435), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_424), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g556 ( .A(n_424), .Y(n_556) );
AND2x2_ASAP7_75t_L g567 ( .A(n_424), .B(n_523), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_424), .B(n_552), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_424), .B(n_554), .Y(n_599) );
AND2x2_ASAP7_75t_L g658 ( .A(n_424), .B(n_603), .Y(n_658) );
INVx4_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g528 ( .A(n_425), .B(n_435), .Y(n_528) );
AND2x2_ASAP7_75t_L g538 ( .A(n_425), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g560 ( .A(n_425), .Y(n_560) );
AND3x2_ASAP7_75t_L g619 ( .A(n_425), .B(n_620), .C(n_621), .Y(n_619) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_435), .Y(n_510) );
INVx1_ASAP7_75t_SL g554 ( .A(n_435), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_435), .B(n_503), .C(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_475), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_445), .A2(n_538), .B(n_590), .C(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_466), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_447), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g606 ( .A(n_447), .Y(n_606) );
AND2x2_ASAP7_75t_L g627 ( .A(n_447), .B(n_477), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_447), .B(n_536), .Y(n_655) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
AND2x2_ASAP7_75t_L g500 ( .A(n_448), .B(n_491), .Y(n_500) );
INVx2_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
AND2x2_ASAP7_75t_L g527 ( .A(n_448), .B(n_477), .Y(n_527) );
AND2x2_ASAP7_75t_L g577 ( .A(n_448), .B(n_466), .Y(n_577) );
INVx1_ASAP7_75t_L g581 ( .A(n_448), .Y(n_581) );
INVx2_ASAP7_75t_SL g491 ( .A(n_457), .Y(n_491) );
BUFx2_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
AND2x2_ASAP7_75t_L g644 ( .A(n_457), .B(n_466), .Y(n_644) );
INVx3_ASAP7_75t_SL g477 ( .A(n_466), .Y(n_477) );
AND2x2_ASAP7_75t_L g499 ( .A(n_466), .B(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g506 ( .A(n_466), .B(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_496), .Y(n_536) );
OR2x2_ASAP7_75t_L g545 ( .A(n_466), .B(n_491), .Y(n_545) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_466), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_521), .Y(n_568) );
AND2x2_ASAP7_75t_L g596 ( .A(n_466), .B(n_479), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_466), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g634 ( .A(n_466), .B(n_478), .Y(n_634) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g558 ( .A(n_477), .B(n_507), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_477), .B(n_500), .Y(n_586) );
AND2x2_ASAP7_75t_L g604 ( .A(n_477), .B(n_521), .Y(n_604) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
AND2x2_ASAP7_75t_L g505 ( .A(n_479), .B(n_491), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_479), .B(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g543 ( .A(n_479), .Y(n_543) );
OR2x2_ASAP7_75t_L g591 ( .A(n_479), .B(n_511), .Y(n_591) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_481), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g497 ( .A(n_483), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_490), .Y(n_498) );
AND2x2_ASAP7_75t_L g526 ( .A(n_491), .B(n_496), .Y(n_526) );
INVx1_ASAP7_75t_L g534 ( .A(n_491), .Y(n_534) );
AND2x2_ASAP7_75t_L g629 ( .A(n_491), .B(n_507), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_501), .B1(n_504), .B2(n_508), .C1(n_512), .C2(n_515), .Y(n_492) );
INVx1_ASAP7_75t_L g624 ( .A(n_493), .Y(n_624) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_499), .Y(n_493) );
AND2x2_ASAP7_75t_L g520 ( .A(n_494), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g531 ( .A(n_494), .B(n_500), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_494), .B(n_522), .Y(n_547) );
OAI222xp33_ASAP7_75t_L g569 ( .A1(n_494), .A2(n_570), .B1(n_575), .B2(n_576), .C1(n_584), .C2(n_586), .Y(n_569) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g557 ( .A(n_496), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_496), .B(n_577), .Y(n_617) );
AND2x2_ASAP7_75t_L g628 ( .A(n_496), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g636 ( .A(n_499), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_501), .B(n_552), .Y(n_615) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_503), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g573 ( .A(n_503), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx3_ASAP7_75t_L g518 ( .A(n_506), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_506), .A2(n_609), .B(n_612), .C(n_614), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_506), .B(n_543), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_506), .B(n_526), .Y(n_648) );
AND2x2_ASAP7_75t_L g521 ( .A(n_507), .B(n_517), .Y(n_521) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g548 ( .A(n_510), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_511), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g600 ( .A(n_511), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g639 ( .A(n_511), .B(n_539), .Y(n_639) );
INVx1_ASAP7_75t_L g651 ( .A(n_511), .Y(n_651) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_514), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g632 ( .A(n_517), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_522), .B(n_524), .C(n_528), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_520), .A2(n_550), .B1(n_565), .B2(n_568), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_521), .B(n_535), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_521), .B(n_543), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_522), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g585 ( .A(n_522), .Y(n_585) );
AND2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_572), .Y(n_592) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
INVxp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NOR4xp25_ASAP7_75t_L g530 ( .A(n_527), .B(n_531), .C(n_532), .D(n_535), .Y(n_530) );
INVx1_ASAP7_75t_SL g601 ( .A(n_528), .Y(n_601) );
AND2x2_ASAP7_75t_L g645 ( .A(n_528), .B(n_646), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_537), .B(n_540), .C(n_549), .Y(n_529) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_536), .B(n_606), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_538), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
INVx1_ASAP7_75t_SL g611 ( .A(n_539), .Y(n_611) );
AND2x2_ASAP7_75t_L g650 ( .A(n_539), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_543), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_547), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_548), .B(n_573), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_555), .B(n_557), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g653 ( .A(n_553), .Y(n_653) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_564), .Y(n_559) );
CKINVDCx16_ASAP7_75t_R g572 ( .A(n_560), .Y(n_572) );
OR2x2_ASAP7_75t_L g610 ( .A(n_560), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g605 ( .A1(n_563), .A2(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_567), .A2(n_594), .B1(n_597), .B2(n_604), .C(n_605), .Y(n_593) );
INVx1_ASAP7_75t_SL g637 ( .A(n_568), .Y(n_637) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OR2x2_ASAP7_75t_L g584 ( .A(n_572), .B(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_L g621 ( .A(n_574), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_581), .B2(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g616 ( .A(n_577), .Y(n_616) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_580), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR4xp25_ASAP7_75t_L g587 ( .A(n_588), .B(n_622), .C(n_635), .D(n_647), .Y(n_587) );
NAND3xp33_ASAP7_75t_SL g588 ( .A(n_589), .B(n_593), .C(n_608), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_591), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_598), .B(n_603), .Y(n_607) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_610), .A2(n_636), .B1(n_637), .B2(n_638), .C(n_640), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_612), .A2(n_627), .B(n_628), .C(n_630), .Y(n_626) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_613), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_630) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_625), .C(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g641 ( .A(n_634), .Y(n_641) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B1(n_652), .B2(n_654), .C(n_656), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g682 ( .A(n_662), .Y(n_682) );
INVx3_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
NAND2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
NOR2xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_SL g693 ( .A(n_673), .Y(n_693) );
INVx1_ASAP7_75t_L g692 ( .A(n_675), .Y(n_692) );
OA21x2_ASAP7_75t_L g695 ( .A1(n_675), .A2(n_693), .B(n_696), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_676), .A2(n_681), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g687 ( .A(n_678), .Y(n_687) );
BUFx2_ASAP7_75t_L g696 ( .A(n_678), .Y(n_696) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
CKINVDCx6p67_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
endmodule