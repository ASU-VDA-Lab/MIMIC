module fake_jpeg_30258_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_6),
.B(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_29),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_86),
.Y(n_114)
);

NOR4xp25_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_60),
.C(n_20),
.D(n_39),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_27),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_49),
.Y(n_86)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_61),
.B1(n_60),
.B2(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_94),
.B1(n_54),
.B2(n_53),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_80),
.B1(n_61),
.B2(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_62),
.B1(n_52),
.B2(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_104),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_67),
.C(n_55),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_114),
.C(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_137)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_54),
.Y(n_104)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_68),
.CON(n_105),
.SN(n_105)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_64),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_0),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_112),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_64),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_3),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_1),
.B(n_2),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_136),
.B(n_120),
.Y(n_143)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_30),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_44),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_38),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_25),
.C(n_31),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_33),
.C(n_36),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_145),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_144),
.C(n_150),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_40),
.CI(n_41),
.CON(n_145),
.SN(n_145)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_43),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_136),
.B1(n_118),
.B2(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_123),
.Y(n_158)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_148),
.A3(n_145),
.B1(n_142),
.B2(n_139),
.C(n_117),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_159),
.B(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_153),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_155),
.B(n_156),
.C(n_151),
.D(n_146),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_122),
.C(n_149),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_121),
.Y(n_165)
);


endmodule