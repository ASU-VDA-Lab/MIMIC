module fake_ariane_2833_n_1097 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_20, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1097);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1097;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_908;
wire n_850;
wire n_788;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_760;
wire n_416;
wire n_969;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_898;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_731;
wire n_336;
wire n_779;
wire n_665;
wire n_903;
wire n_754;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_821;
wire n_561;
wire n_928;
wire n_770;
wire n_839;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_894;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_538;
wire n_352;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_543;
wire n_362;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_774;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_115),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_150),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_48),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_114),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_170),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_257),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_18),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_135),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_187),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_255),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_9),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_47),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_112),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_57),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_75),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_146),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_74),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_103),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_122),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_100),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_13),
.Y(n_318)
);

BUFx2_ASAP7_75t_SL g319 ( 
.A(n_106),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_147),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_154),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_142),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_5),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_263),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_40),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_210),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_246),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_174),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_212),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_127),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_13),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_73),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_140),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_196),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_131),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_157),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_177),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_151),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_78),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_232),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_207),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_3),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_275),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_70),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_2),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_211),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_277),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_134),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_23),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_32),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_240),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_133),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_205),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_225),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_19),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_105),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_197),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_267),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_82),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_102),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_273),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_162),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_34),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_92),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_14),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_178),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_42),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_1),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_259),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_49),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_172),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_117),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_124),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_31),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_233),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_279),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_130),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_23),
.Y(n_386)
);

CKINVDCx12_ASAP7_75t_R g387 ( 
.A(n_90),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_282),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_271),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_76),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_280),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_143),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_182),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_60),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_107),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_18),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_61),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_116),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_238),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_272),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_164),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_17),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_269),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_46),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_113),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_229),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_208),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_168),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_149),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_185),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_141),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_118),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_4),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_128),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_71),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_87),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_190),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_123),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_2),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_260),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_200),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_50),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_8),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_4),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_91),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_67),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_226),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_137),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_244),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_15),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_192),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_53),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_95),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_30),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_223),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_9),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_8),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_22),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_25),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_63),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_62),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_43),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_125),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_241),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_108),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_268),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_222),
.Y(n_448)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_55),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_27),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_11),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_256),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_179),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_94),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_217),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_262),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_204),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_274),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_126),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_261),
.Y(n_460)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_158),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_230),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_88),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_41),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_39),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_51),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_44),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_248),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_121),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_167),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_236),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_144),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_258),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_281),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_342),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_357),
.B(n_0),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_357),
.B(n_0),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_360),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_374),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_324),
.B(n_1),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_292),
.B(n_3),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_342),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_293),
.B(n_6),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_7),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_297),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_290),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_306),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_358),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_326),
.B(n_7),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_303),
.B(n_10),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_358),
.B(n_10),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_322),
.B(n_33),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_303),
.B(n_11),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_345),
.B(n_12),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_301),
.B(n_12),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_290),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_298),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_320),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_345),
.B(n_14),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_308),
.B(n_15),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_333),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_392),
.B(n_406),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_290),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_381),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_323),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_381),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_347),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_309),
.B(n_16),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_310),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_381),
.Y(n_523)
);

BUFx8_ASAP7_75t_SL g524 ( 
.A(n_440),
.Y(n_524)
);

BUFx8_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_314),
.B(n_16),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_318),
.B(n_19),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_444),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_321),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_304),
.B(n_20),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_327),
.B(n_20),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_429),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_328),
.B(n_21),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_338),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_344),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_350),
.B(n_356),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_361),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_307),
.B(n_21),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_365),
.B(n_22),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_349),
.B(n_24),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_367),
.B(n_24),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_354),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

BUFx8_ASAP7_75t_SL g545 ( 
.A(n_341),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_311),
.B(n_25),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_346),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_355),
.B(n_26),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_335),
.B(n_26),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_336),
.B(n_27),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_368),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_337),
.B(n_364),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_371),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_375),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_376),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_377),
.B(n_28),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_351),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_394),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_409),
.B(n_28),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_378),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_289),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_379),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_388),
.B(n_29),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_390),
.B(n_29),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_397),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_382),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_386),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_396),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_401),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_403),
.B(n_405),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_413),
.B(n_30),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_422),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_458),
.B(n_35),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_412),
.B(n_415),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_387),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_31),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_428),
.B(n_32),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_435),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_434),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_441),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_483),
.A2(n_456),
.B1(n_468),
.B2(n_446),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_479),
.A2(n_438),
.B1(n_439),
.B2(n_437),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_476),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_478),
.A2(n_474),
.B1(n_451),
.B2(n_450),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_510),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_480),
.A2(n_366),
.B1(n_414),
.B2(n_448),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_481),
.A2(n_454),
.B1(n_457),
.B2(n_455),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_495),
.A2(n_467),
.B1(n_469),
.B2(n_460),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_492),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_493),
.B(n_319),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_470),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_545),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_291),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_561),
.B(n_472),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_477),
.A2(n_473),
.B1(n_471),
.B2(n_466),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_294),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

AO22x2_ASAP7_75t_L g599 ( 
.A1(n_496),
.A2(n_449),
.B1(n_461),
.B2(n_463),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_498),
.A2(n_465),
.B1(n_464),
.B2(n_462),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_475),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_500),
.A2(n_461),
.B1(n_449),
.B2(n_453),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_482),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_482),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_491),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_494),
.A2(n_373),
.B1(n_459),
.B2(n_452),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_540),
.A2(n_370),
.B1(n_296),
.B2(n_445),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_489),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_295),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_548),
.A2(n_572),
.B1(n_511),
.B2(n_501),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_299),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_520),
.A2(n_380),
.B1(n_302),
.B2(n_443),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_503),
.B(n_300),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_506),
.B(n_305),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_513),
.B(n_312),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_497),
.A2(n_449),
.B1(n_461),
.B2(n_442),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_489),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_527),
.A2(n_575),
.B1(n_571),
.B2(n_505),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_514),
.A2(n_383),
.B1(n_315),
.B2(n_436),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_SL g620 ( 
.A1(n_487),
.A2(n_384),
.B1(n_316),
.B2(n_433),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_513),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_547),
.A2(n_372),
.B1(n_317),
.B2(n_432),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_513),
.B(n_313),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_553),
.A2(n_385),
.B1(n_325),
.B2(n_427),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_530),
.A2(n_389),
.B1(n_329),
.B2(n_421),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_530),
.A2(n_369),
.B1(n_330),
.B2(n_418),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_538),
.A2(n_449),
.B1(n_461),
.B2(n_417),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_547),
.A2(n_363),
.B1(n_331),
.B2(n_416),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_538),
.A2(n_549),
.B1(n_550),
.B2(n_546),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_573),
.A2(n_391),
.B1(n_332),
.B2(n_411),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_490),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_576),
.B(n_334),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_546),
.A2(n_393),
.B1(n_340),
.B2(n_410),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_512),
.A2(n_556),
.B1(n_564),
.B2(n_577),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_518),
.B(n_339),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_543),
.B(n_343),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_576),
.B(n_348),
.Y(n_638)
);

OAI22xp33_ASAP7_75t_L g639 ( 
.A1(n_573),
.A2(n_399),
.B1(n_353),
.B2(n_408),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_549),
.A2(n_400),
.B1(n_359),
.B2(n_407),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_550),
.A2(n_559),
.B1(n_579),
.B2(n_569),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_509),
.B(n_352),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_559),
.A2(n_404),
.B1(n_395),
.B2(n_362),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_485),
.A2(n_461),
.B1(n_449),
.B2(n_38),
.Y(n_644)
);

OAI22xp33_ASAP7_75t_L g645 ( 
.A1(n_566),
.A2(n_461),
.B1(n_449),
.B2(n_45),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_552),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_646)
);

AO22x2_ASAP7_75t_L g647 ( 
.A1(n_552),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_647)
);

AND2x2_ASAP7_75t_SL g648 ( 
.A(n_531),
.B(n_59),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_502),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_521),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_570),
.B(n_69),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_526),
.A2(n_563),
.B1(n_539),
.B2(n_555),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_555),
.A2(n_72),
.B1(n_77),
.B2(n_79),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_SL g654 ( 
.A1(n_533),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_568),
.B(n_84),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_515),
.B(n_85),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_605),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_582),
.B(n_528),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_R g659 ( 
.A(n_593),
.B(n_515),
.Y(n_659)
);

INVx3_ASAP7_75t_R g660 ( 
.A(n_584),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_649),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_601),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_607),
.B(n_522),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_629),
.B(n_534),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_591),
.B(n_606),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_586),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_599),
.B(n_557),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_535),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_634),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_610),
.B(n_537),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_598),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_603),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_641),
.B(n_504),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_551),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_621),
.B(n_519),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_618),
.B(n_522),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_604),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_608),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_581),
.B(n_529),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_554),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_636),
.Y(n_683)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_599),
.B(n_524),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_617),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_590),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_636),
.B(n_542),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_596),
.B(n_560),
.Y(n_689)
);

XOR2xp5_ASAP7_75t_L g690 ( 
.A(n_602),
.B(n_646),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_590),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_635),
.B(n_558),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_656),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_632),
.B(n_504),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_595),
.B(n_536),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_580),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_588),
.B(n_614),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g698 ( 
.A(n_602),
.B(n_562),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_592),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_651),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_637),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_594),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_597),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_611),
.B(n_507),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_638),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_655),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_646),
.Y(n_709)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_637),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_647),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_613),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_647),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_616),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_644),
.Y(n_715)
);

AND2x6_ASAP7_75t_L g716 ( 
.A(n_625),
.B(n_507),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_614),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_615),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_616),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_R g721 ( 
.A(n_623),
.B(n_578),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_612),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_654),
.Y(n_724)
);

XNOR2x2_ASAP7_75t_L g725 ( 
.A(n_626),
.B(n_525),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_633),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_640),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_643),
.B(n_562),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_624),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_619),
.B(n_558),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_583),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_600),
.B(n_558),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_622),
.B(n_567),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_653),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_628),
.Y(n_737)
);

AND2x4_ASAP7_75t_SL g738 ( 
.A(n_717),
.B(n_674),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_695),
.B(n_565),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_680),
.B(n_630),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_704),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_704),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_639),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_671),
.B(n_565),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_664),
.B(n_609),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_661),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_677),
.B(n_484),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_694),
.B(n_677),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_679),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_696),
.A2(n_650),
.B(n_488),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_675),
.B(n_567),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_670),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_687),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_709),
.B(n_574),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_659),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_708),
.B(n_574),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_712),
.B(n_525),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_683),
.B(n_574),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_706),
.B(n_508),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_672),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_699),
.A2(n_541),
.B(n_532),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_674),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_673),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_666),
.B(n_516),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_703),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_692),
.A2(n_541),
.B(n_532),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_728),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_516),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_685),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_724),
.B(n_519),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_689),
.B(n_517),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_658),
.B(n_517),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_523),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_686),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_724),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_723),
.B(n_523),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_718),
.B(n_544),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_681),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_711),
.B(n_544),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_726),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_702),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_713),
.B(n_86),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_716),
.B(n_519),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_669),
.B(n_532),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_705),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_710),
.B(n_541),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_729),
.B(n_89),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_692),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_707),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_727),
.B(n_93),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_691),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_732),
.B(n_96),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_720),
.B(n_97),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_737),
.B(n_98),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_724),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_716),
.B(n_288),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

BUFx4f_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_693),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_736),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_700),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_719),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_734),
.B(n_99),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_716),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_698),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_731),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_730),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_730),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_779),
.Y(n_813)
);

INVx6_ASAP7_75t_L g814 ( 
.A(n_779),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_806),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_740),
.B(n_665),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_779),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_768),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_779),
.B(n_697),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_804),
.B(n_690),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_738),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_757),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_744),
.B(n_722),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_738),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_765),
.B(n_701),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_786),
.B(n_735),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_772),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_745),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_784),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_769),
.A2(n_733),
.B(n_735),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_806),
.Y(n_831)
);

NAND2x1_ASAP7_75t_L g832 ( 
.A(n_799),
.B(n_676),
.Y(n_832)
);

INVx5_ASAP7_75t_L g833 ( 
.A(n_799),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_804),
.B(n_733),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_739),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_807),
.B(n_676),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_789),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_772),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_807),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_772),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_801),
.B(n_662),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_801),
.B(n_725),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_745),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_785),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_767),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_763),
.A2(n_721),
.B(n_668),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_768),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_740),
.B(n_684),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_742),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_804),
.B(n_688),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_776),
.Y(n_851)
);

NAND2x1_ASAP7_75t_SL g852 ( 
.A(n_807),
.B(n_688),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_749),
.B(n_799),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_742),
.B(n_660),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_764),
.B(n_101),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_743),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_768),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_747),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_750),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_743),
.B(n_104),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_817),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_817),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_822),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_824),
.Y(n_864)
);

BUFx2_ASAP7_75t_R g865 ( 
.A(n_846),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_827),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_817),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_817),
.Y(n_868)
);

BUFx2_ASAP7_75t_SL g869 ( 
.A(n_821),
.Y(n_869)
);

INVx5_ASAP7_75t_L g870 ( 
.A(n_814),
.Y(n_870)
);

INVx6_ASAP7_75t_L g871 ( 
.A(n_833),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_814),
.Y(n_872)
);

INVx5_ASAP7_75t_L g873 ( 
.A(n_814),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_816),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_858),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_833),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_826),
.A2(n_786),
.B1(n_746),
.B2(n_741),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_815),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_833),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_831),
.Y(n_880)
);

CKINVDCx14_ASAP7_75t_R g881 ( 
.A(n_825),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_859),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_837),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_833),
.Y(n_884)
);

BUFx4f_ASAP7_75t_SL g885 ( 
.A(n_844),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_839),
.B(n_813),
.Y(n_886)
);

BUFx4_ASAP7_75t_SL g887 ( 
.A(n_854),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_854),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_839),
.B(n_748),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_838),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_841),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_813),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_887),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_877),
.A2(n_826),
.B1(n_823),
.B2(n_848),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_889),
.A2(n_823),
.B1(n_846),
.B2(n_812),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_885),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_889),
.B(n_811),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_888),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_878),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_875),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_883),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_879),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_881),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_863),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_881),
.B(n_829),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_874),
.A2(n_791),
.B1(n_830),
.B2(n_794),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_882),
.Y(n_907)
);

INVx8_ASAP7_75t_L g908 ( 
.A(n_870),
.Y(n_908)
);

INVx6_ASAP7_75t_L g909 ( 
.A(n_870),
.Y(n_909)
);

OAI22xp33_ASAP7_75t_L g910 ( 
.A1(n_874),
.A2(n_850),
.B1(n_842),
.B2(n_853),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_SL g911 ( 
.A1(n_891),
.A2(n_850),
.B(n_751),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_876),
.Y(n_912)
);

OAI22xp33_ASAP7_75t_L g913 ( 
.A1(n_891),
.A2(n_842),
.B1(n_853),
.B2(n_843),
.Y(n_913)
);

AND2x4_ASAP7_75t_SL g914 ( 
.A(n_872),
.B(n_841),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_882),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_880),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_892),
.A2(n_829),
.B1(n_843),
.B2(n_792),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_SL g918 ( 
.A1(n_865),
.A2(n_842),
.B1(n_820),
.B2(n_830),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_866),
.A2(n_834),
.B1(n_805),
.B2(n_803),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_880),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_905),
.B(n_866),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_903),
.B(n_890),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_896),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_894),
.A2(n_906),
.B1(n_895),
.B2(n_910),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_906),
.A2(n_791),
.B1(n_794),
.B2(n_798),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_894),
.A2(n_917),
.B1(n_897),
.B2(n_911),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_918),
.A2(n_809),
.B1(n_820),
.B2(n_845),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_SL g928 ( 
.A1(n_893),
.A2(n_895),
.B1(n_904),
.B2(n_852),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_898),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_899),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_912),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_900),
.B(n_890),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_901),
.B(n_849),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_910),
.A2(n_798),
.B1(n_771),
.B2(n_828),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_914),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_914),
.B(n_849),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_913),
.A2(n_834),
.B1(n_796),
.B2(n_797),
.Y(n_937)
);

OAI22xp33_ASAP7_75t_L g938 ( 
.A1(n_913),
.A2(n_805),
.B1(n_803),
.B2(n_739),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_919),
.A2(n_836),
.B1(n_810),
.B2(n_851),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_912),
.B(n_864),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_919),
.A2(n_808),
.B1(n_836),
.B2(n_886),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_908),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_916),
.A2(n_810),
.B1(n_783),
.B2(n_753),
.Y(n_943)
);

INVx4_ASAP7_75t_SL g944 ( 
.A(n_909),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_920),
.B(n_748),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_909),
.A2(n_886),
.B1(n_796),
.B2(n_797),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_908),
.Y(n_947)
);

AOI222xp33_ASAP7_75t_L g948 ( 
.A1(n_907),
.A2(n_840),
.B1(n_783),
.B2(n_756),
.C1(n_775),
.C2(n_752),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_907),
.A2(n_819),
.B1(n_759),
.B2(n_739),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_902),
.A2(n_856),
.B1(n_800),
.B2(n_841),
.Y(n_950)
);

OAI221xp5_ASAP7_75t_L g951 ( 
.A1(n_925),
.A2(n_781),
.B1(n_790),
.B2(n_864),
.C(n_856),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_946),
.A2(n_781),
.B(n_855),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_932),
.B(n_912),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_926),
.B(n_912),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_924),
.A2(n_802),
.B1(n_778),
.B2(n_754),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_924),
.A2(n_802),
.B1(n_754),
.B2(n_773),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_928),
.A2(n_773),
.B1(n_770),
.B2(n_774),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_930),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_927),
.A2(n_770),
.B1(n_774),
.B2(n_915),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_948),
.A2(n_770),
.B1(n_795),
.B2(n_886),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_937),
.A2(n_770),
.B1(n_795),
.B2(n_886),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_950),
.A2(n_886),
.B1(n_756),
.B2(n_869),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_934),
.A2(n_766),
.B1(n_762),
.B2(n_755),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_SL g964 ( 
.A1(n_936),
.A2(n_760),
.B1(n_909),
.B2(n_908),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_938),
.A2(n_755),
.B1(n_857),
.B2(n_847),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_938),
.A2(n_818),
.B1(n_835),
.B2(n_780),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_943),
.A2(n_835),
.B1(n_793),
.B2(n_860),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_949),
.A2(n_793),
.B1(n_777),
.B2(n_761),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_SL g969 ( 
.A1(n_921),
.A2(n_760),
.B1(n_758),
.B2(n_787),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_939),
.A2(n_761),
.B1(n_758),
.B2(n_788),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_945),
.A2(n_761),
.B1(n_832),
.B2(n_854),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_940),
.B(n_892),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_923),
.A2(n_892),
.B1(n_902),
.B2(n_871),
.Y(n_973)
);

OAI22xp33_ASAP7_75t_L g974 ( 
.A1(n_941),
.A2(n_870),
.B1(n_873),
.B2(n_879),
.Y(n_974)
);

OAI221xp5_ASAP7_75t_L g975 ( 
.A1(n_933),
.A2(n_782),
.B1(n_861),
.B2(n_867),
.C(n_872),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_931),
.B(n_861),
.Y(n_976)
);

OAI222xp33_ASAP7_75t_L g977 ( 
.A1(n_935),
.A2(n_861),
.B1(n_867),
.B2(n_879),
.C1(n_884),
.C2(n_870),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_947),
.A2(n_867),
.B1(n_884),
.B2(n_870),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_884),
.B1(n_873),
.B2(n_862),
.Y(n_979)
);

AOI221xp5_ASAP7_75t_L g980 ( 
.A1(n_929),
.A2(n_942),
.B1(n_868),
.B2(n_862),
.C(n_873),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_954),
.B(n_944),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_954),
.B(n_944),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_953),
.B(n_944),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_SL g984 ( 
.A1(n_951),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.C(n_120),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_972),
.B(n_862),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_972),
.B(n_862),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_974),
.B(n_868),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_952),
.A2(n_873),
.B(n_868),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_975),
.B(n_873),
.C(n_868),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_976),
.B(n_979),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_287),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_973),
.B(n_129),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_980),
.B(n_132),
.C(n_136),
.Y(n_993)
);

XOR2xp5_ASAP7_75t_L g994 ( 
.A(n_978),
.B(n_286),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_L g995 ( 
.A1(n_957),
.A2(n_138),
.B(n_139),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_961),
.B(n_145),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_958),
.B(n_285),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_962),
.B(n_148),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_SL g999 ( 
.A1(n_977),
.A2(n_152),
.B(n_153),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_955),
.B(n_283),
.Y(n_1000)
);

AOI211xp5_ASAP7_75t_L g1001 ( 
.A1(n_969),
.A2(n_155),
.B(n_156),
.C(n_159),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_964),
.B(n_161),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_971),
.B(n_163),
.C(n_165),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_956),
.B(n_166),
.C(n_169),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_960),
.A2(n_171),
.B1(n_173),
.B2(n_176),
.Y(n_1005)
);

OAI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_963),
.A2(n_181),
.B(n_183),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_984),
.B(n_966),
.C(n_967),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_986),
.Y(n_1008)
);

OAI211xp5_ASAP7_75t_SL g1009 ( 
.A1(n_991),
.A2(n_959),
.B(n_970),
.C(n_965),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_985),
.B(n_968),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_990),
.B(n_184),
.Y(n_1011)
);

INVxp33_ASAP7_75t_SL g1012 ( 
.A(n_983),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_981),
.Y(n_1013)
);

AOI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_998),
.A2(n_1006),
.B1(n_996),
.B2(n_999),
.C(n_989),
.Y(n_1014)
);

NAND4xp75_ASAP7_75t_L g1015 ( 
.A(n_1002),
.B(n_186),
.C(n_188),
.D(n_189),
.Y(n_1015)
);

OA211x2_ASAP7_75t_L g1016 ( 
.A1(n_1002),
.A2(n_191),
.B(n_193),
.C(n_194),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_1001),
.B(n_198),
.C(n_199),
.Y(n_1017)
);

NAND4xp75_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_202),
.C(n_203),
.D(n_206),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_982),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_987),
.B(n_988),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_987),
.B(n_209),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_992),
.B(n_213),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_1012),
.B(n_994),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1008),
.B(n_997),
.Y(n_1024)
);

NAND4xp75_ASAP7_75t_L g1025 ( 
.A(n_1014),
.B(n_1000),
.C(n_995),
.D(n_996),
.Y(n_1025)
);

XOR2x2_ASAP7_75t_L g1026 ( 
.A(n_1007),
.B(n_1003),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_993),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1013),
.B(n_1022),
.Y(n_1028)
);

XOR2x2_ASAP7_75t_L g1029 ( 
.A(n_1007),
.B(n_1004),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1020),
.B(n_1005),
.Y(n_1030)
);

NAND4xp75_ASAP7_75t_L g1031 ( 
.A(n_1016),
.B(n_214),
.C(n_215),
.D(n_216),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_278),
.Y(n_1032)
);

INVxp67_ASAP7_75t_SL g1033 ( 
.A(n_1010),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_218),
.Y(n_1034)
);

XOR2x2_ASAP7_75t_L g1035 ( 
.A(n_1017),
.B(n_219),
.Y(n_1035)
);

XNOR2xp5_ASAP7_75t_L g1036 ( 
.A(n_1018),
.B(n_220),
.Y(n_1036)
);

XNOR2xp5_ASAP7_75t_L g1037 ( 
.A(n_1015),
.B(n_221),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1021),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_1024),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_1027),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1038),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1033),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1027),
.Y(n_1043)
);

XNOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1030),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1029),
.A2(n_224),
.B1(n_227),
.B2(n_231),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_1032),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1032),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_1028),
.Y(n_1049)
);

XNOR2x2_ASAP7_75t_L g1050 ( 
.A(n_1025),
.B(n_234),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1023),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1034),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1044),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

AO22x1_ASAP7_75t_L g1055 ( 
.A1(n_1040),
.A2(n_1035),
.B1(n_1036),
.B2(n_1037),
.Y(n_1055)
);

OA22x2_ASAP7_75t_L g1056 ( 
.A1(n_1040),
.A2(n_1031),
.B1(n_239),
.B2(n_243),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_1039),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_1052),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_1047),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1041),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1048),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1043),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1045),
.A2(n_235),
.B1(n_245),
.B2(n_247),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_1049),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1048),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1043),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_SL g1068 ( 
.A(n_1053),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1061),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1063),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1067),
.Y(n_1072)
);

AOI22x1_ASAP7_75t_L g1073 ( 
.A1(n_1069),
.A2(n_1061),
.B1(n_1053),
.B2(n_1067),
.Y(n_1073)
);

AOI221x1_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_1054),
.B1(n_1066),
.B2(n_1058),
.C(n_1062),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_1071),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1072),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1068),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1076),
.Y(n_1078)
);

OA22x2_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_1065),
.B1(n_1068),
.B2(n_1059),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1075),
.A2(n_1045),
.B1(n_1056),
.B2(n_1055),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1080),
.B(n_1059),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1078),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1079),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1081),
.B(n_1058),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1082),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1084),
.Y(n_1087)
);

AO22x2_ASAP7_75t_L g1088 ( 
.A1(n_1087),
.A2(n_1083),
.B1(n_1074),
.B2(n_1073),
.Y(n_1088)
);

INVxp67_ASAP7_75t_SL g1089 ( 
.A(n_1088),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_1085),
.B1(n_1086),
.B2(n_1056),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1090),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_1050),
.B1(n_1047),
.B2(n_1060),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1093),
.A2(n_1064),
.B1(n_1046),
.B2(n_1057),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

AOI221xp5_ASAP7_75t_L g1096 ( 
.A1(n_1095),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.C(n_254),
.Y(n_1096)
);

AOI211xp5_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_264),
.B(n_265),
.C(n_266),
.Y(n_1097)
);


endmodule