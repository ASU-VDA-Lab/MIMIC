module fake_jpeg_24283_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_7),
.B(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_6),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_24),
.Y(n_90)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_42),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_85),
.B1(n_86),
.B2(n_92),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_18),
.B1(n_30),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_24),
.B1(n_37),
.B2(n_25),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_69),
.Y(n_104)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_18),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_87),
.B1(n_43),
.B2(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_91),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_43),
.B1(n_47),
.B2(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_18),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_49),
.B1(n_56),
.B2(n_37),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_126),
.B1(n_72),
.B2(n_84),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_43),
.B1(n_64),
.B2(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_112),
.B1(n_118),
.B2(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_53),
.C(n_39),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_121),
.C(n_93),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_53),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_116),
.B(n_93),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_65),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_128),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_64),
.B1(n_61),
.B2(n_65),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_79),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_44),
.B(n_49),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_120),
.B1(n_127),
.B2(n_67),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_39),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_39),
.B1(n_48),
.B2(n_47),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_25),
.B1(n_22),
.B2(n_26),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_44),
.Y(n_128)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_130),
.Y(n_184)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_0),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_143),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_156),
.B1(n_118),
.B2(n_112),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_145),
.Y(n_172)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_34),
.B(n_22),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_152),
.B1(n_119),
.B2(n_108),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_106),
.B(n_121),
.Y(n_162)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_86),
.B1(n_34),
.B2(n_26),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_38),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_40),
.B1(n_46),
.B2(n_45),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_173),
.B1(n_176),
.B2(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_159),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_165),
.B(n_174),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_121),
.B(n_115),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_117),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_31),
.C(n_21),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_100),
.B1(n_79),
.B2(n_60),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_40),
.B1(n_107),
.B2(n_114),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_40),
.B1(n_114),
.B2(n_108),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_40),
.B1(n_95),
.B2(n_69),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_154),
.B(n_136),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_132),
.A3(n_156),
.B1(n_135),
.B2(n_143),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_149),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_40),
.B1(n_92),
.B2(n_46),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_38),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_94),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_28),
.B1(n_36),
.B2(n_45),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_142),
.B1(n_141),
.B2(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_45),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_74),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_38),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_213),
.B(n_160),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_184),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_192),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_144),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_196),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_38),
.A3(n_46),
.B1(n_48),
.B2(n_47),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_205),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_202),
.B1(n_47),
.B2(n_48),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_28),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_31),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_8),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_200),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_31),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_7),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_204),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_20),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_83),
.C(n_48),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_32),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_16),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_21),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_219),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_0),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_0),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_16),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_158),
.B(n_16),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_1),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_21),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_31),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_201),
.C(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_233),
.C(n_192),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_171),
.B1(n_173),
.B2(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_179),
.B1(n_169),
.B2(n_159),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_208),
.B1(n_195),
.B2(n_194),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_176),
.C(n_164),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_166),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_238),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_187),
.B(n_1),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_242),
.B(n_217),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_32),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_217),
.B1(n_195),
.B2(n_111),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_33),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_13),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_246),
.A2(n_247),
.B1(n_238),
.B2(n_33),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_250),
.B1(n_253),
.B2(n_256),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_212),
.B(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_238),
.C(n_230),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_199),
.B1(n_197),
.B2(n_111),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_71),
.B1(n_47),
.B2(n_33),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_227),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_31),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_244),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_33),
.C(n_32),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_241),
.C(n_239),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_221),
.B1(n_233),
.B2(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_222),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_271),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_222),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_221),
.B1(n_226),
.B2(n_229),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_276),
.B1(n_284),
.B2(n_262),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_253),
.B(n_246),
.C(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_231),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_282),
.C(n_260),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_231),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_32),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_290),
.Y(n_302)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_255),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_1),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_291),
.C(n_294),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_273),
.C(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_259),
.C(n_265),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_27),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_303),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_297),
.B(n_270),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_309),
.C(n_310),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_27),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_299),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_294),
.C(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_320),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_285),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_296),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_296),
.C(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_285),
.B1(n_298),
.B2(n_1),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_4),
.Y(n_331)
);

OAI322xp33_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_10),
.Y(n_324)
);

AO22x1_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_4),
.B1(n_10),
.B2(n_12),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_313),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_3),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_23),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_322),
.A3(n_330),
.B1(n_326),
.B2(n_321),
.C1(n_27),
.C2(n_23),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_322),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_10),
.C(n_12),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_23),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_27),
.Y(n_339)
);


endmodule