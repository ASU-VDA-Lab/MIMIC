module fake_jpeg_2641_n_126 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_17),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_55),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_38),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_41),
.Y(n_71)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2x1p5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_60),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_91),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_42),
.B(n_34),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_2),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_0),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_70),
.C(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_105),
.B1(n_5),
.B2(n_10),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_4),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_27),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_30),
.B(n_31),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_21),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_28),
.B1(n_6),
.B2(n_8),
.C(n_9),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_5),
.B(n_13),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_114),
.C(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_102),
.C(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_112),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_119),
.B(n_107),
.C(n_112),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_108),
.B(n_115),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule