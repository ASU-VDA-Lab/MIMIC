module fake_jpeg_1646_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_55),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_50),
.B1(n_45),
.B2(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_73),
.B1(n_57),
.B2(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_54),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_38),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_63),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_52),
.B1(n_47),
.B2(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_61),
.B1(n_56),
.B2(n_66),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_80),
.B1(n_79),
.B2(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_73),
.B1(n_71),
.B2(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_55),
.B(n_66),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_48),
.B(n_42),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_59),
.B1(n_52),
.B2(n_61),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_59),
.B1(n_56),
.B2(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_105),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_103),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_46),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_0),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_118),
.B(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_0),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_35),
.B1(n_32),
.B2(n_30),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_17),
.B(n_34),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_48),
.B1(n_42),
.B2(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_29),
.C(n_26),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_120),
.C(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_25),
.B(n_24),
.C(n_23),
.D(n_21),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_20),
.B(n_19),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_123),
.C(n_132),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_104),
.B1(n_6),
.B2(n_8),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_125),
.B1(n_126),
.B2(n_8),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_132),
.B1(n_134),
.B2(n_123),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_147),
.B(n_139),
.C(n_141),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_148),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_135),
.B1(n_131),
.B2(n_126),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_140),
.C(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_147),
.Y(n_153)
);

AOI31xp33_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_153),
.A3(n_149),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_139),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_143),
.B(n_6),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_5),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_5),
.A3(n_9),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_155),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_14),
.Y(n_159)
);


endmodule