module fake_jpeg_6078_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_14),
.B1(n_24),
.B2(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_19),
.B1(n_24),
.B2(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_40),
.B1(n_44),
.B2(n_15),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_50),
.B1(n_13),
.B2(n_55),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_28),
.B(n_27),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_27),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_30),
.B(n_28),
.C(n_45),
.D(n_31),
.Y(n_62)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_34),
.B1(n_45),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_68),
.B1(n_56),
.B2(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_57),
.B1(n_50),
.B2(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_34),
.B1(n_32),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_48),
.B1(n_34),
.B2(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_89),
.B1(n_27),
.B2(n_21),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_84),
.B1(n_65),
.B2(n_74),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_51),
.B1(n_32),
.B2(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_12),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_31),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_60),
.C(n_62),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_60),
.B(n_72),
.C(n_27),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_21),
.B1(n_9),
.B2(n_11),
.Y(n_99)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_86),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_78),
.B(n_76),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_100),
.C(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_93),
.A3(n_85),
.B1(n_82),
.B2(n_76),
.C1(n_94),
.C2(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.C(n_116),
.Y(n_120)
);

OAI321xp33_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_100),
.A3(n_97),
.B1(n_77),
.B2(n_79),
.C(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_25),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_104),
.B1(n_110),
.B2(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_105),
.C(n_108),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_105),
.C(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_7),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_23),
.Y(n_126)
);

OAI221xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_2),
.C(n_3),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_23),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_10),
.C(n_3),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_4),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_125),
.C(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_128),
.Y(n_137)
);


endmodule