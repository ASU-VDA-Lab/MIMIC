module fake_jpeg_4694_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_60),
.B1(n_64),
.B2(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_24),
.B1(n_32),
.B2(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_56),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_26),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_69),
.Y(n_77)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_95),
.B1(n_99),
.B2(n_15),
.Y(n_125)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_33),
.B1(n_22),
.B2(n_43),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_23),
.B1(n_25),
.B2(n_2),
.Y(n_127)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_17),
.B1(n_54),
.B2(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_84),
.B(n_98),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_31),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_35),
.B1(n_28),
.B2(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_17),
.B1(n_65),
.B2(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_0),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_27),
.B(n_38),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_73),
.B(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_72),
.B1(n_57),
.B2(n_65),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_114),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_97),
.B(n_82),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_57),
.B1(n_67),
.B2(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_110),
.B1(n_111),
.B2(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_113),
.B1(n_116),
.B2(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_77),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_70),
.B1(n_51),
.B2(n_67),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_25),
.Y(n_152)
);

AOI22x1_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_43),
.B1(n_54),
.B2(n_38),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_33),
.B1(n_22),
.B2(n_46),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_90),
.B1(n_86),
.B2(n_84),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_33),
.A3(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_88),
.B(n_77),
.C(n_89),
.D(n_25),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_76),
.B1(n_79),
.B2(n_88),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_127),
.B1(n_78),
.B2(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_95),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_138),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_158),
.B(n_114),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_85),
.B1(n_95),
.B2(n_89),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_127),
.B(n_121),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_92),
.C(n_96),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_151),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_156),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_110),
.B1(n_105),
.B2(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_94),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_113),
.B1(n_127),
.B2(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_88),
.C(n_89),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_0),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_0),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_1),
.C(n_2),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_1),
.B(n_2),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_151),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_152),
.CI(n_184),
.CON(n_204),
.SN(n_204)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_181),
.B(n_185),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_184),
.B1(n_154),
.B2(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_131),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_124),
.B1(n_125),
.B2(n_111),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_187),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_140),
.B1(n_135),
.B2(n_151),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_197),
.B1(n_203),
.B2(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_150),
.B1(n_136),
.B2(n_117),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_202),
.B1(n_209),
.B2(n_167),
.Y(n_231)
);

XNOR2x2_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_198),
.B(n_204),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_145),
.B1(n_140),
.B2(n_133),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_158),
.B(n_137),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_137),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_205),
.C(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_101),
.B1(n_139),
.B2(n_154),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_152),
.C(n_109),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_156),
.B(n_155),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_163),
.A2(n_107),
.B1(n_108),
.B2(n_122),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_129),
.B1(n_123),
.B2(n_130),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_159),
.B1(n_169),
.B2(n_175),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_217),
.B(n_218),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_181),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_219),
.B(n_231),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_213),
.B1(n_209),
.B2(n_179),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_220),
.Y(n_253)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_205),
.C(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_228),
.B(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_237),
.Y(n_260)
);

OAI22x1_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_178),
.B1(n_160),
.B2(n_186),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_234),
.B1(n_130),
.B2(n_123),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_160),
.B1(n_187),
.B2(n_170),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_166),
.B1(n_159),
.B2(n_164),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_236),
.B1(n_192),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_182),
.B1(n_169),
.B2(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_123),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_257),
.CI(n_225),
.CON(n_279),
.SN(n_279)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_192),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_256),
.B(n_245),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_248),
.C(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_200),
.C(n_191),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_177),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_190),
.C(n_177),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_171),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_201),
.C(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_256),
.C(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_201),
.C(n_166),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_216),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_228),
.B1(n_236),
.B2(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_1),
.C(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_219),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_260),
.B(n_251),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_218),
.B1(n_232),
.B2(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_240),
.B1(n_242),
.B2(n_230),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_275),
.B1(n_276),
.B2(n_282),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_234),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_277),
.B(n_279),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_264),
.B(n_257),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_280),
.B(n_284),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_246),
.A2(n_223),
.B(n_241),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_5),
.C(n_6),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_252),
.C(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_14),
.B(n_7),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_249),
.C(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_263),
.C(n_6),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_278),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_12),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_268),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_304),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_266),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_278),
.C(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_279),
.Y(n_309)
);

NAND2x1_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_267),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_311),
.B1(n_11),
.B2(n_7),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_279),
.B1(n_283),
.B2(n_282),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_287),
.B1(n_298),
.B2(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_318),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_5),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_5),
.B(n_7),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_311),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_11),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_325),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_328),
.C(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_305),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_310),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_332),
.C(n_11),
.Y(n_337)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_321),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_8),
.B(n_9),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_306),
.B1(n_9),
.B2(n_11),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.C(n_327),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_334),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_335),
.B(n_333),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_8),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_8),
.B(n_9),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_8),
.Y(n_344)
);


endmodule