module fake_jpeg_23661_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx2_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_54),
.Y(n_90)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_27),
.B2(n_20),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_71),
.B1(n_32),
.B2(n_19),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_35),
.B1(n_33),
.B2(n_27),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_74),
.B1(n_84),
.B2(n_23),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_35),
.B1(n_27),
.B2(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_25),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_17),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_34),
.B1(n_18),
.B2(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_38),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_17),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_29),
.B1(n_24),
.B2(n_37),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_95),
.B1(n_10),
.B2(n_15),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_26),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_103),
.B(n_25),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_52),
.B(n_37),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_2),
.C(n_4),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_77),
.B(n_81),
.C(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_34),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_48),
.A3(n_37),
.B1(n_51),
.B2(n_49),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_30),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_37),
.B1(n_32),
.B2(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_109),
.B1(n_110),
.B2(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_106),
.Y(n_137)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_37),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_37),
.B1(n_23),
.B2(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_72),
.B1(n_55),
.B2(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_113),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_62),
.B(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_115),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_31),
.B1(n_19),
.B2(n_28),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_28),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_63),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_83),
.B1(n_79),
.B2(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_139),
.B1(n_157),
.B2(n_129),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_131),
.B(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_128),
.B(n_141),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_134),
.B1(n_150),
.B2(n_111),
.Y(n_186)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_136),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_1),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_60),
.B(n_67),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_109),
.B1(n_97),
.B2(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_63),
.B1(n_30),
.B2(n_4),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_14),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_9),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_144),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_90),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_90),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_106),
.B1(n_117),
.B2(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_119),
.Y(n_191)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_10),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_154),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_8),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_100),
.C(n_88),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_95),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_148),
.B(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_174),
.B1(n_186),
.B2(n_157),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_91),
.B(n_92),
.C(n_90),
.D(n_87),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_181),
.C(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_168),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_92),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_171),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_140),
.B(n_124),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_88),
.B1(n_92),
.B2(n_109),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_173),
.B1(n_144),
.B2(n_130),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_98),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_123),
.A2(n_109),
.B1(n_108),
.B2(n_111),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_131),
.Y(n_208)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_137),
.Y(n_189)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_141),
.B(n_125),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_199),
.B(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_198),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_133),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_136),
.B1(n_139),
.B2(n_128),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_213),
.B1(n_216),
.B2(n_220),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_212),
.B(n_215),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_146),
.B(n_125),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_131),
.B(n_145),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_210),
.B(n_164),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_171),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_134),
.B1(n_119),
.B2(n_101),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_214),
.B1(n_160),
.B2(n_176),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_178),
.B(n_169),
.Y(n_210)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_135),
.B1(n_120),
.B2(n_107),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_101),
.B1(n_149),
.B2(n_107),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_170),
.A2(n_89),
.B1(n_135),
.B2(n_5),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_162),
.A2(n_5),
.B(n_7),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_7),
.B1(n_12),
.B2(n_14),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_228),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_173),
.B1(n_185),
.B2(n_175),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_231),
.B1(n_237),
.B2(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_159),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_167),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_238),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_193),
.A2(n_201),
.B1(n_200),
.B2(n_198),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_236),
.B(n_220),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_211),
.B1(n_212),
.B2(n_195),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_246),
.B1(n_247),
.B2(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_207),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_210),
.B1(n_192),
.B2(n_222),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_221),
.B1(n_194),
.B2(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_231),
.B1(n_225),
.B2(n_224),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_197),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_260),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_199),
.C(n_203),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_265),
.C(n_165),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_208),
.B1(n_205),
.B2(n_168),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_267),
.B1(n_228),
.B2(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_203),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_262),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_177),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_217),
.B1(n_163),
.B2(n_188),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_263),
.B(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_163),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_218),
.B1(n_161),
.B2(n_190),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_179),
.B1(n_165),
.B2(n_7),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_238),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_277),
.C(n_281),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_243),
.B(n_242),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_280),
.B(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_274),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_276),
.B1(n_248),
.B2(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_226),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_223),
.B1(n_246),
.B2(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_232),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_283),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_232),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_285),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_246),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_165),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_251),
.C(n_261),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_298),
.C(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_282),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_299),
.B(n_269),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_254),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_259),
.C(n_250),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_281),
.C(n_282),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_308),
.B(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_274),
.CI(n_272),
.CON(n_305),
.SN(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_294),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_309),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_276),
.C(n_284),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_179),
.B1(n_255),
.B2(n_15),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.C(n_300),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_295),
.B1(n_286),
.B2(n_289),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_319),
.B(n_322),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_311),
.A2(n_304),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_321),
.B(n_303),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_326)
);

OAI31xp33_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_312),
.A3(n_314),
.B(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_301),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_315),
.B(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_326),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_315),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_307),
.B1(n_15),
.B2(n_16),
.Y(n_332)
);


endmodule