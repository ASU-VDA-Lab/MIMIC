module real_aes_1333_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g563 ( .A(n_0), .B(n_218), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_1), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g141 ( .A(n_2), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_3), .B(n_500), .Y(n_499) );
NAND2xp33_ASAP7_75t_SL g555 ( .A(n_4), .B(n_158), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_5), .B(n_202), .Y(n_210) );
INVx1_ASAP7_75t_L g548 ( .A(n_6), .Y(n_548) );
INVx1_ASAP7_75t_L g149 ( .A(n_7), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g834 ( .A(n_8), .Y(n_834) );
OAI22x1_ASAP7_75t_R g793 ( .A1(n_9), .A2(n_77), .B1(n_794), .B2(n_795), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_9), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_10), .Y(n_175) );
AND2x2_ASAP7_75t_L g497 ( .A(n_11), .B(n_190), .Y(n_497) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g219 ( .A(n_14), .Y(n_219) );
AOI221x1_ASAP7_75t_L g551 ( .A1(n_15), .A2(n_162), .B1(n_502), .B2(n_552), .C(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_16), .B(n_500), .Y(n_535) );
INVx1_ASAP7_75t_L g117 ( .A(n_17), .Y(n_117) );
INVx1_ASAP7_75t_L g216 ( .A(n_18), .Y(n_216) );
INVx1_ASAP7_75t_SL g231 ( .A(n_19), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_20), .B(n_152), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_21), .A2(n_27), .B1(n_488), .B2(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_21), .Y(n_824) );
AOI33xp33_ASAP7_75t_L g256 ( .A1(n_22), .A2(n_51), .A3(n_136), .B1(n_144), .B2(n_257), .B3(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_23), .A2(n_502), .B(n_503), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_24), .B(n_218), .Y(n_504) );
AOI221xp5_ASAP7_75t_SL g527 ( .A1(n_25), .A2(n_41), .B1(n_500), .B2(n_502), .C(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g167 ( .A(n_26), .Y(n_167) );
NOR3xp33_ASAP7_75t_L g120 ( .A(n_27), .B(n_121), .C(n_312), .Y(n_120) );
INVx1_ASAP7_75t_SL g488 ( .A(n_27), .Y(n_488) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_28), .A2(n_90), .B(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g191 ( .A(n_28), .B(n_90), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_29), .B(n_221), .Y(n_539) );
INVxp67_ASAP7_75t_L g550 ( .A(n_30), .Y(n_550) );
AND2x2_ASAP7_75t_L g523 ( .A(n_31), .B(n_189), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_32), .B(n_142), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_33), .A2(n_502), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_34), .B(n_221), .Y(n_529) );
INVx1_ASAP7_75t_L g135 ( .A(n_35), .Y(n_135) );
AND2x2_ASAP7_75t_L g147 ( .A(n_35), .B(n_138), .Y(n_147) );
AND2x2_ASAP7_75t_L g158 ( .A(n_35), .B(n_141), .Y(n_158) );
OR2x6_ASAP7_75t_L g115 ( .A(n_36), .B(n_116), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g832 ( .A(n_36), .B(n_833), .C(n_835), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_37), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_38), .B(n_142), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_39), .A2(n_163), .B1(n_198), .B2(n_202), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_40), .B(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_42), .A2(n_81), .B1(n_133), .B2(n_502), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_43), .B(n_152), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_44), .B(n_218), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_45), .B(n_129), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_46), .B(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_47), .Y(n_201) );
AND2x2_ASAP7_75t_L g566 ( .A(n_48), .B(n_189), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_49), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_50), .B(n_189), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_52), .B(n_152), .Y(n_187) );
INVx1_ASAP7_75t_L g140 ( .A(n_53), .Y(n_140) );
INVx1_ASAP7_75t_L g154 ( .A(n_53), .Y(n_154) );
AND2x2_ASAP7_75t_L g188 ( .A(n_54), .B(n_189), .Y(n_188) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_55), .A2(n_73), .B1(n_133), .B2(n_142), .C(n_148), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_56), .B(n_142), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_57), .B(n_500), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_58), .B(n_163), .Y(n_177) );
AOI21xp5_ASAP7_75t_SL g240 ( .A1(n_59), .A2(n_133), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g514 ( .A(n_60), .B(n_189), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_61), .B(n_221), .Y(n_564) );
INVx1_ASAP7_75t_L g213 ( .A(n_62), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_63), .B(n_218), .Y(n_512) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_64), .B(n_190), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_65), .A2(n_502), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g186 ( .A(n_66), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_67), .B(n_221), .Y(n_505) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_68), .B(n_129), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_69), .A2(n_133), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g138 ( .A(n_70), .Y(n_138) );
INVx1_ASAP7_75t_L g156 ( .A(n_70), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_71), .B(n_142), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_72), .A2(n_103), .B1(n_829), .B2(n_837), .Y(n_102) );
AND2x2_ASAP7_75t_L g233 ( .A(n_74), .B(n_162), .Y(n_233) );
INVx1_ASAP7_75t_L g214 ( .A(n_75), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_76), .A2(n_133), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_77), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_78), .A2(n_133), .B(n_204), .C(n_208), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_79), .B(n_500), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_80), .A2(n_84), .B1(n_142), .B2(n_500), .Y(n_576) );
INVx1_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_82), .B(n_117), .Y(n_836) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_83), .B(n_162), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_85), .A2(n_133), .B1(n_254), .B2(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_86), .B(n_218), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_87), .B(n_218), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_88), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_89), .A2(n_502), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g242 ( .A(n_91), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_92), .B(n_221), .Y(n_511) );
AND2x2_ASAP7_75t_L g260 ( .A(n_93), .B(n_162), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_94), .A2(n_165), .B(n_166), .C(n_169), .Y(n_164) );
INVxp67_ASAP7_75t_L g553 ( .A(n_95), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_96), .B(n_500), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_97), .B(n_221), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_98), .A2(n_502), .B(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_SL g106 ( .A(n_99), .Y(n_106) );
BUFx2_ASAP7_75t_L g809 ( .A(n_99), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_100), .B(n_152), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g821 ( .A1(n_101), .A2(n_822), .B1(n_823), .B2(n_825), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_101), .Y(n_822) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B(n_806), .Y(n_103) );
CKINVDCx11_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx8_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_801), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_792), .B(n_796), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_119), .B1(n_490), .B2(n_788), .Y(n_109) );
CKINVDCx6p67_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_111), .Y(n_805) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
AND2x6_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g790 ( .A(n_114), .B(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_L g800 ( .A(n_114), .B(n_115), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_114), .B(n_791), .Y(n_815) );
CKINVDCx16_ASAP7_75t_R g835 ( .A(n_114), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_115), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AOI211xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_383), .B(n_486), .C(n_489), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_120), .A2(n_383), .B(n_486), .Y(n_803) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_122), .A2(n_384), .B(n_488), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g819 ( .A(n_122), .B(n_461), .Y(n_819) );
NOR2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_290), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_273), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_192), .B1(n_234), .B2(n_248), .C(n_263), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_179), .Y(n_125) );
NAND2x1_ASAP7_75t_SL g299 ( .A(n_126), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g326 ( .A(n_126), .B(n_296), .Y(n_326) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_126), .Y(n_372) );
AND2x2_ASAP7_75t_L g380 ( .A(n_126), .B(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g484 ( .A(n_126), .Y(n_484) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_160), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_128), .Y(n_262) );
INVx1_ASAP7_75t_L g278 ( .A(n_128), .Y(n_278) );
AND2x4_ASAP7_75t_L g285 ( .A(n_128), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_128), .B(n_160), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_128), .B(n_281), .Y(n_322) );
INVx1_ASAP7_75t_L g333 ( .A(n_128), .Y(n_333) );
INVxp67_ASAP7_75t_L g367 ( .A(n_128), .Y(n_367) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_159), .Y(n_128) );
INVx2_ASAP7_75t_SL g208 ( .A(n_129), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_129), .A2(n_535), .B(n_536), .Y(n_534) );
BUFx4f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_131), .B(n_191), .Y(n_190) );
AND2x4_ASAP7_75t_L g202 ( .A(n_131), .B(n_191), .Y(n_202) );
INVxp67_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_133), .A2(n_142), .B1(n_547), .B2(n_549), .Y(n_546) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
NOR2x1p5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
INVx1_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x6_ASAP7_75t_L g150 ( .A(n_137), .B(n_144), .Y(n_150) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g218 ( .A(n_138), .B(n_153), .Y(n_218) );
AND2x6_ASAP7_75t_L g502 ( .A(n_139), .B(n_147), .Y(n_502) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx2_ASAP7_75t_L g144 ( .A(n_140), .Y(n_144) );
AND2x4_ASAP7_75t_L g221 ( .A(n_140), .B(n_155), .Y(n_221) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_141), .Y(n_145) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_146), .Y(n_142) );
INVx1_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVxp33_ASAP7_75t_L g257 ( .A(n_144), .Y(n_257) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_150), .B(n_151), .C(n_157), .Y(n_148) );
INVxp67_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_150), .A2(n_157), .B(n_186), .C(n_187), .Y(n_185) );
INVx2_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_150), .A2(n_168), .B1(n_213), .B2(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_150), .A2(n_157), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_150), .A2(n_157), .B(n_242), .C(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
AND2x4_ASAP7_75t_L g500 ( .A(n_152), .B(n_158), .Y(n_500) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_157), .A2(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_157), .B(n_202), .Y(n_222) );
INVx1_ASAP7_75t_L g254 ( .A(n_157), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_157), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_157), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_157), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_157), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_157), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_157), .A2(n_563), .B(n_564), .Y(n_562) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_158), .Y(n_169) );
INVx2_ASAP7_75t_L g250 ( .A(n_160), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_160), .B(n_181), .Y(n_266) );
INVx1_ASAP7_75t_L g284 ( .A(n_160), .Y(n_284) );
INVx1_ASAP7_75t_L g331 ( .A(n_160), .Y(n_331) );
OR2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_172), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B1(n_170), .B2(n_171), .Y(n_161) );
INVx3_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_163), .B(n_174), .Y(n_173) );
AOI21x1_ASAP7_75t_L g559 ( .A1(n_163), .A2(n_560), .B(n_566), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_168), .B(n_202), .C(n_555), .Y(n_554) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_171), .A2(n_182), .B(n_188), .Y(n_181) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_171), .A2(n_182), .B(n_188), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_179), .B(n_303), .Y(n_308) );
AND2x2_ASAP7_75t_L g320 ( .A(n_179), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g339 ( .A(n_179), .B(n_285), .Y(n_339) );
INVx1_ASAP7_75t_L g348 ( .A(n_179), .Y(n_348) );
AND2x2_ASAP7_75t_L g396 ( .A(n_179), .B(n_295), .Y(n_396) );
OR2x2_ASAP7_75t_L g439 ( .A(n_179), .B(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x4_ASAP7_75t_L g279 ( .A(n_180), .B(n_280), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_180), .B(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g261 ( .A(n_181), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_181), .B(n_281), .Y(n_359) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_181), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_189), .Y(n_226) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_189), .A2(n_527), .B(n_531), .Y(n_526) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_223), .Y(n_193) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_194), .B(n_318), .Y(n_363) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g325 ( .A(n_195), .B(n_316), .Y(n_325) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_209), .Y(n_195) );
INVx1_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
AND2x4_ASAP7_75t_L g271 ( .A(n_196), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_196), .Y(n_311) );
AND2x2_ASAP7_75t_L g481 ( .A(n_196), .B(n_237), .Y(n_481) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_203), .Y(n_196) );
NOR3xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .C(n_201), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_202), .A2(n_240), .B(n_244), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_202), .A2(n_499), .B(n_501), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_202), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_202), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_202), .B(n_553), .Y(n_552) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_208), .A2(n_252), .B(n_260), .Y(n_251) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_208), .A2(n_252), .B(n_260), .Y(n_281) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_208), .A2(n_575), .B(n_578), .Y(n_574) );
INVx3_ASAP7_75t_L g272 ( .A(n_209), .Y(n_272) );
INVx2_ASAP7_75t_L g289 ( .A(n_209), .Y(n_289) );
NOR2x1_ASAP7_75t_SL g306 ( .A(n_209), .B(n_237), .Y(n_306) );
AND2x2_ASAP7_75t_L g344 ( .A(n_209), .B(n_225), .Y(n_344) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_215), .B(n_222), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B1(n_219), .B2(n_220), .Y(n_215) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g418 ( .A(n_223), .Y(n_418) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g247 ( .A(n_224), .Y(n_247) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
INVx1_ASAP7_75t_L g316 ( .A(n_225), .Y(n_316) );
INVx1_ASAP7_75t_L g376 ( .A(n_225), .Y(n_376) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_225), .Y(n_395) );
OR2x2_ASAP7_75t_L g401 ( .A(n_225), .B(n_237), .Y(n_401) );
AND2x2_ASAP7_75t_L g445 ( .A(n_225), .B(n_272), .Y(n_445) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_233), .Y(n_225) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_226), .A2(n_508), .B(n_514), .Y(n_507) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_226), .A2(n_517), .B(n_523), .Y(n_516) );
AO21x2_ASAP7_75t_L g655 ( .A1(n_226), .A2(n_517), .B(n_523), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_246), .Y(n_235) );
AND2x2_ASAP7_75t_L g287 ( .A(n_236), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g441 ( .A(n_236), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g446 ( .A(n_236), .Y(n_446) );
AND2x2_ASAP7_75t_L g458 ( .A(n_236), .B(n_344), .Y(n_458) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_245), .Y(n_236) );
INVx4_ASAP7_75t_L g269 ( .A(n_237), .Y(n_269) );
INVx2_ASAP7_75t_L g319 ( .A(n_237), .Y(n_319) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_237), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_237), .B(n_377), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_237), .B(n_247), .Y(n_450) );
AND2x2_ASAP7_75t_L g476 ( .A(n_237), .B(n_289), .Y(n_476) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x4_ASAP7_75t_L g378 ( .A(n_245), .B(n_269), .Y(n_378) );
AND2x2_ASAP7_75t_L g305 ( .A(n_246), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_246), .B(n_310), .Y(n_323) );
INVx1_ASAP7_75t_L g357 ( .A(n_246), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_246), .B(n_271), .Y(n_413) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_247), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_248), .A2(n_330), .B1(n_474), .B2(n_477), .Y(n_473) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_261), .Y(n_248) );
INVx1_ASAP7_75t_L g403 ( .A(n_249), .Y(n_403) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g277 ( .A(n_250), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g426 ( .A(n_250), .B(n_298), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_250), .B(n_298), .Y(n_435) );
INVx2_ASAP7_75t_L g286 ( .A(n_251), .Y(n_286) );
AND2x4_ASAP7_75t_L g296 ( .A(n_251), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_251), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_253), .B(n_259), .Y(n_252) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_262), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_265), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g370 ( .A(n_265), .B(n_285), .Y(n_370) );
INVx2_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g408 ( .A(n_266), .B(n_322), .Y(n_408) );
INVxp33_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g389 ( .A(n_268), .Y(n_389) );
NOR2x1_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_269), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_269), .Y(n_335) );
INVx2_ASAP7_75t_L g399 ( .A(n_270), .Y(n_399) );
NAND2xp33_ASAP7_75t_SL g474 ( .A(n_270), .B(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g340 ( .A(n_271), .B(n_319), .Y(n_340) );
AND2x2_ASAP7_75t_L g274 ( .A(n_272), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g377 ( .A(n_272), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B1(n_282), .B2(n_287), .Y(n_273) );
AND2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g407 ( .A(n_274), .Y(n_407) );
INVx1_ASAP7_75t_L g356 ( .A(n_275), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_276), .A2(n_315), .B1(n_320), .B2(n_323), .Y(n_314) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx2_ASAP7_75t_L g440 ( .A(n_277), .Y(n_440) );
BUFx3_ASAP7_75t_L g405 ( .A(n_278), .Y(n_405) );
INVx1_ASAP7_75t_L g428 ( .A(n_279), .Y(n_428) );
AND2x2_ASAP7_75t_L g366 ( .A(n_280), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g433 ( .A(n_280), .B(n_298), .Y(n_433) );
INVx1_ASAP7_75t_L g467 ( .A(n_280), .Y(n_467) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI21xp33_ASAP7_75t_L g304 ( .A1(n_282), .A2(n_305), .B(n_307), .Y(n_304) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_282), .A2(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g415 ( .A(n_284), .Y(n_415) );
AND2x2_ASAP7_75t_L g432 ( .A(n_284), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g422 ( .A(n_285), .B(n_381), .Y(n_422) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g434 ( .A(n_285), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g379 ( .A(n_288), .B(n_378), .Y(n_379) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_289), .B(n_318), .Y(n_317) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_289), .B(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_301), .B(n_304), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_299), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_294), .A2(n_310), .B1(n_335), .B2(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_298), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_300), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_300), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g442 ( .A(n_303), .Y(n_442) );
AND2x2_ASAP7_75t_L g429 ( .A(n_306), .B(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_R g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_310), .B(n_393), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_312), .Y(n_487) );
OR3x2_ASAP7_75t_L g818 ( .A(n_312), .B(n_385), .C(n_819), .Y(n_818) );
NAND3x1_ASAP7_75t_SL g312 ( .A(n_313), .B(n_327), .C(n_341), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_324), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_315), .A2(n_425), .B1(n_427), .B2(n_429), .Y(n_424) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_316), .B(n_355), .Y(n_369) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_321), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g390 ( .A(n_321), .B(n_331), .Y(n_390) );
AND2x2_ASAP7_75t_L g414 ( .A(n_321), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_325), .A2(n_421), .B(n_422), .Y(n_420) );
AND2x2_ASAP7_75t_L g472 ( .A(n_325), .B(n_351), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_326), .A2(n_479), .B1(n_482), .B2(n_485), .Y(n_478) );
AOI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_334), .B(n_338), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
BUFx2_ASAP7_75t_L g448 ( .A(n_331), .Y(n_448) );
INVx1_ASAP7_75t_SL g455 ( .A(n_331), .Y(n_455) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_332), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_361), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B(n_349), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_344), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_344), .B(n_355), .Y(n_436) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_352), .B(n_358), .Y(n_349) );
OR2x6_ASAP7_75t_L g406 ( .A(n_351), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g456 ( .A(n_359), .Y(n_456) );
OR2x2_ASAP7_75t_L g483 ( .A(n_359), .B(n_484), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_360), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_371), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_368), .B2(n_370), .Y(n_362) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_365), .Y(n_463) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_379), .B2(n_380), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
AND2x4_ASAP7_75t_SL g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_459), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_409), .C(n_437), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_397), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_391), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp33_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_402), .B1(n_406), .B2(n_408), .Y(n_397) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_399), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_401), .B(n_407), .Y(n_477) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx3_ASAP7_75t_L g465 ( .A(n_405), .Y(n_465) );
INVx2_ASAP7_75t_L g469 ( .A(n_406), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_423), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_420), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_419), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_424), .B(n_431), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_426), .B(n_467), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g451 ( .A(n_434), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B(n_443), .C(n_452), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g470 ( .A1(n_440), .A2(n_471), .B(n_473), .C(n_478), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B1(n_449), .B2(n_451), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_459), .A2(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_462), .B(n_470), .Y(n_461) );
AOI21xp33_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B(n_468), .Y(n_462) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_489), .B(n_805), .Y(n_804) );
AO22x2_ASAP7_75t_L g802 ( .A1(n_490), .A2(n_789), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_699), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_621), .C(n_671), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_588), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_524), .B1(n_541), .B2(n_571), .C(n_580), .Y(n_494) );
INVx1_ASAP7_75t_SL g670 ( .A(n_495), .Y(n_670) );
AND2x4_ASAP7_75t_SL g495 ( .A(n_496), .B(n_506), .Y(n_495) );
INVx2_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
OR2x2_ASAP7_75t_L g614 ( .A(n_496), .B(n_605), .Y(n_614) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_496), .Y(n_629) );
INVx5_ASAP7_75t_L g636 ( .A(n_496), .Y(n_636) );
AND2x4_ASAP7_75t_L g642 ( .A(n_496), .B(n_516), .Y(n_642) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_496), .B(n_573), .Y(n_645) );
OR2x2_ASAP7_75t_L g654 ( .A(n_496), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g661 ( .A(n_496), .B(n_507), .Y(n_661) );
AND2x2_ASAP7_75t_L g762 ( .A(n_496), .B(n_515), .Y(n_762) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx3_ASAP7_75t_SL g613 ( .A(n_506), .Y(n_613) );
AND2x2_ASAP7_75t_L g657 ( .A(n_506), .B(n_573), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_506), .A2(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g698 ( .A(n_506), .B(n_636), .Y(n_698) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_507), .B(n_516), .Y(n_579) );
OR2x2_ASAP7_75t_L g583 ( .A(n_507), .B(n_516), .Y(n_583) );
INVx1_ASAP7_75t_L g591 ( .A(n_507), .Y(n_591) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_507), .Y(n_603) );
INVx2_ASAP7_75t_L g611 ( .A(n_507), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_507), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g720 ( .A(n_507), .B(n_605), .Y(n_720) );
AND2x2_ASAP7_75t_L g735 ( .A(n_507), .B(n_573), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_513), .Y(n_508) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g604 ( .A(n_516), .B(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_516), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_524), .B(n_728), .Y(n_727) );
NOR2x1p5_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g557 ( .A(n_526), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_526), .B(n_533), .Y(n_586) );
INVx1_ASAP7_75t_L g596 ( .A(n_526), .Y(n_596) );
INVx2_ASAP7_75t_L g619 ( .A(n_526), .Y(n_619) );
INVx2_ASAP7_75t_L g625 ( .A(n_526), .Y(n_625) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_526), .Y(n_695) );
OR2x2_ASAP7_75t_L g726 ( .A(n_526), .B(n_533), .Y(n_726) );
OR2x2_ASAP7_75t_L g742 ( .A(n_532), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_SL g544 ( .A(n_533), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g569 ( .A(n_533), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g606 ( .A(n_533), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g618 ( .A(n_533), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g631 ( .A(n_533), .B(n_597), .Y(n_631) );
OR2x2_ASAP7_75t_L g639 ( .A(n_533), .B(n_545), .Y(n_639) );
INVx2_ASAP7_75t_L g666 ( .A(n_533), .Y(n_666) );
INVx1_ASAP7_75t_L g684 ( .A(n_533), .Y(n_684) );
NOR2xp33_ASAP7_75t_R g717 ( .A(n_533), .B(n_558), .Y(n_717) );
OR2x6_ASAP7_75t_L g533 ( .A(n_534), .B(n_540), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_567), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_542), .A2(n_609), .B1(n_612), .B2(n_615), .Y(n_608) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_556), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g623 ( .A(n_544), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g658 ( .A(n_544), .B(n_659), .Y(n_658) );
AND2x4_ASAP7_75t_L g737 ( .A(n_544), .B(n_715), .Y(n_737) );
INVx3_ASAP7_75t_L g570 ( .A(n_545), .Y(n_570) );
AND2x4_ASAP7_75t_L g597 ( .A(n_545), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_545), .B(n_558), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_545), .B(n_619), .Y(n_664) );
AND2x2_ASAP7_75t_L g669 ( .A(n_545), .B(n_666), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_545), .B(n_557), .Y(n_706) );
INVx1_ASAP7_75t_L g776 ( .A(n_545), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_545), .B(n_694), .Y(n_787) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g568 ( .A(n_558), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_558), .B(n_570), .Y(n_587) );
INVx2_ASAP7_75t_L g598 ( .A(n_558), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_558), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g640 ( .A(n_558), .B(n_619), .Y(n_640) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_558), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_558), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g729 ( .A(n_558), .Y(n_729) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_568), .B(n_596), .Y(n_607) );
AOI221x1_ASAP7_75t_SL g701 ( .A1(n_569), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_711), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_569), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g759 ( .A(n_569), .B(n_624), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_569), .B(n_781), .Y(n_780) );
OR2x2_ASAP7_75t_L g690 ( .A(n_570), .B(n_618), .Y(n_690) );
AND2x2_ASAP7_75t_L g728 ( .A(n_570), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_579), .Y(n_572) );
AND2x2_ASAP7_75t_L g581 ( .A(n_573), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g676 ( .A(n_573), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_573), .B(n_592), .Y(n_681) );
AND2x4_ASAP7_75t_L g710 ( .A(n_573), .B(n_611), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_573), .B(n_642), .Y(n_746) );
OR2x2_ASAP7_75t_L g764 ( .A(n_573), .B(n_695), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_573), .B(n_655), .Y(n_774) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g605 ( .A(n_574), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g630 ( .A(n_579), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_579), .A2(n_638), .B1(n_641), .B2(n_643), .Y(n_637) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx2_ASAP7_75t_L g593 ( .A(n_581), .Y(n_593) );
AND2x2_ASAP7_75t_L g732 ( .A(n_582), .B(n_592), .Y(n_732) );
AND2x2_ASAP7_75t_L g778 ( .A(n_582), .B(n_645), .Y(n_778) );
AND2x2_ASAP7_75t_L g783 ( .A(n_582), .B(n_634), .Y(n_783) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI32xp33_ASAP7_75t_L g752 ( .A1(n_584), .A2(n_654), .A3(n_734), .B1(n_753), .B2(n_755), .Y(n_752) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
AOI211xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_594), .B(n_599), .C(n_608), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_593), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_591), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_592), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g772 ( .A(n_592), .Y(n_772) );
AND2x2_ASAP7_75t_L g682 ( .A(n_594), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_SL g594 ( .A(n_595), .B(n_597), .Y(n_594) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_595), .Y(n_782) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_596), .Y(n_651) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_596), .Y(n_751) );
INVx1_ASAP7_75t_L g648 ( .A(n_597), .Y(n_648) );
AND2x2_ASAP7_75t_L g714 ( .A(n_597), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_597), .B(n_725), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_601), .A2(n_681), .B(n_682), .Y(n_680) );
AND2x2_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g610 ( .A(n_605), .B(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g634 ( .A(n_605), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_610), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g741 ( .A(n_610), .Y(n_741) );
AND2x2_ASAP7_75t_L g771 ( .A(n_610), .B(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_611), .Y(n_748) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_613), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g688 ( .A(n_614), .Y(n_688) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g647 ( .A(n_618), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_619), .Y(n_715) );
AND2x2_ASAP7_75t_L g724 ( .A(n_620), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_644), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_631), .B2(n_632), .C(n_637), .Y(n_622) );
INVx1_ASAP7_75t_L g743 ( .A(n_624), .Y(n_743) );
INVxp33_ASAP7_75t_SL g775 ( .A(n_624), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_626), .A2(n_722), .B(n_730), .Y(n_721) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_630), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g643 ( .A(n_631), .Y(n_643) );
AND2x2_ASAP7_75t_L g678 ( .A(n_631), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_631), .A2(n_759), .B1(n_760), .B2(n_763), .Y(n_758) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
OR2x2_ASAP7_75t_L g653 ( .A(n_634), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_634), .B(n_642), .Y(n_692) );
AND2x4_ASAP7_75t_L g709 ( .A(n_636), .B(n_655), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_636), .B(n_710), .Y(n_756) );
AND2x2_ASAP7_75t_L g768 ( .A(n_636), .B(n_720), .Y(n_768) );
NAND2xp33_ASAP7_75t_L g753 ( .A(n_638), .B(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_SL g696 ( .A(n_639), .Y(n_696) );
INVx1_ASAP7_75t_L g767 ( .A(n_640), .Y(n_767) );
INVx2_ASAP7_75t_SL g719 ( .A(n_642), .Y(n_719) );
AOI211xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B(n_649), .C(n_667), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B(n_656), .C(n_660), .Y(n_649) );
OR2x6_ASAP7_75t_SL g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g679 ( .A(n_651), .Y(n_679) );
INVx1_ASAP7_75t_SL g704 ( .A(n_654), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_654), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_659), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g745 ( .A1(n_663), .A2(n_746), .B1(n_747), .B2(n_749), .Y(n_745) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_677), .B(n_680), .C(n_685), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_691), .B2(n_693), .C(n_697), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g777 ( .A1(n_696), .A2(n_778), .B1(n_779), .B2(n_783), .C1(n_784), .C2(n_786), .Y(n_777) );
INVx2_ASAP7_75t_L g712 ( .A(n_698), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_738), .C(n_757), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_721), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_709), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_710), .B(n_772), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_716), .B2(n_718), .Y(n_711) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVxp33_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_719), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_727), .A2(n_731), .B1(n_733), .B2(n_736), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_742), .B(n_744), .C(n_752), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_765), .C(n_777), .Y(n_757) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_769), .B(n_776), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_773), .B(n_775), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVxp33_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_793), .B(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B(n_826), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_816), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
BUFx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx2_ASAP7_75t_L g828 ( .A(n_815), .Y(n_828) );
AOI22x1_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_820), .B2(n_821), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g825 ( .A(n_823), .Y(n_825) );
INVx1_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
BUFx8_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
BUFx4f_ASAP7_75t_SL g838 ( .A(n_831), .Y(n_838) );
NAND2xp5_ASAP7_75t_SL g831 ( .A(n_832), .B(n_836), .Y(n_831) );
BUFx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
endmodule