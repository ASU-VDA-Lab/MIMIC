module fake_netlist_5_451_n_2124 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2124);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2124;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2009;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_1079;
wire n_457;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_101),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_73),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_62),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_76),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_103),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_159),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_30),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_78),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_108),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_133),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_32),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_171),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_86),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_63),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_141),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_35),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_69),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_194),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_175),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_2),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_74),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_23),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_119),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_88),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_36),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_32),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_117),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_57),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_123),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_59),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_184),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_112),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_62),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_90),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_116),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_102),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_92),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_87),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_89),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_33),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_82),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_150),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_163),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_109),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_8),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_149),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_114),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_162),
.Y(n_291)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_144),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_57),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_35),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_121),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_65),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_75),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_173),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_37),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_95),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_3),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_8),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_160),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_29),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_193),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_45),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_66),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_51),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_135),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_157),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_13),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_25),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_132),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_26),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_4),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_28),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_45),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_93),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_31),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_110),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_111),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_30),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_10),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_151),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_139),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_36),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_142),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_44),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_14),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_48),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_12),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_18),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_127),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_113),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_67),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_66),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_131),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_10),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_26),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_21),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_204),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_42),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_15),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_71),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_100),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_49),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_50),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_77),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_61),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_60),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_59),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_24),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_11),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_27),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_180),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_99),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_197),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_168),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_13),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_165),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_181),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_70),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_155),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_39),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_84),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_50),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_152),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_20),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_14),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_128),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_49),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_200),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_83),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_12),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_192),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_33),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_154),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_107),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_146),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_5),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_6),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_64),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_125),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_105),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_72),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_40),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_196),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_147),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_18),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_46),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_42),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_80),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_167),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_183),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_136),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_34),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_44),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_138),
.Y(n_410)
);

BUFx8_ASAP7_75t_SL g411 ( 
.A(n_96),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_364),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_225),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_281),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_281),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_411),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_281),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_281),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_281),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_233),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_246),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_310),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_310),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_303),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_250),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_310),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_304),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_244),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_310),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_310),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_331),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_299),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_251),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_309),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_252),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_256),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_339),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_253),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_209),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_219),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_318),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_313),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_215),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_275),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_240),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_245),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_351),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_261),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_320),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_248),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_276),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_406),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_271),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_272),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_287),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_290),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_294),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_280),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_305),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_253),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_307),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_213),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_264),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_312),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_330),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_228),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_327),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_273),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_332),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_340),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_348),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_282),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_289),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_352),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_366),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_273),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_285),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_273),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_259),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_231),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_259),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_218),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_213),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_253),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_288),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_291),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_218),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_293),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_258),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_210),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_268),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_298),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_316),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_268),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_407),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_231),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_273),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_296),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_328),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_416),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_429),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_436),
.B(n_375),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_391),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_497),
.B(n_231),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_443),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_445),
.B(n_224),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_368),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_412),
.A2(n_314),
.B1(n_409),
.B2(n_224),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_476),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_418),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_421),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_446),
.B(n_404),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_476),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_456),
.Y(n_544)
);

NOR2x1_ASAP7_75t_L g545 ( 
.A(n_499),
.B(n_368),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_507),
.B(n_368),
.Y(n_546)
);

BUFx6f_ASAP7_75t_SL g547 ( 
.A(n_463),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_419),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_420),
.B(n_375),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_435),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_446),
.B(n_248),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_464),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_424),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_424),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_384),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_471),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_430),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_430),
.B(n_384),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_207),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_431),
.B(n_207),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_448),
.B(n_248),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_433),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_492),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_214),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_448),
.B(n_255),
.C(n_243),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_434),
.B(n_208),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_438),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_450),
.B(n_249),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_439),
.B(n_440),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_481),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_499),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_508),
.A2(n_344),
.B(n_296),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_508),
.B(n_344),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_489),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_511),
.B(n_367),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_489),
.A2(n_377),
.B(n_367),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_425),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_428),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_515),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_450),
.B(n_208),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_503),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_573),
.B(n_505),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_598),
.B(n_509),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_582),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_524),
.B(n_414),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_524),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_523),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_563),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_506),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_527),
.B(n_510),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_518),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_528),
.B(n_531),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_522),
.B(n_516),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_543),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

AND3x2_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_397),
.C(n_377),
.Y(n_616)
);

INVx6_ASAP7_75t_L g617 ( 
.A(n_521),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_528),
.B(n_452),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_529),
.B(n_473),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_519),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_520),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_548),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_548),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_547),
.B(n_486),
.Y(n_628)
);

NOR2x1p5_ASAP7_75t_L g629 ( 
.A(n_544),
.B(n_417),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_532),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_534),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_564),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_555),
.B(n_473),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_534),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_538),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

BUFx6f_ASAP7_75t_SL g638 ( 
.A(n_523),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_527),
.B(n_264),
.Y(n_639)
);

AND2x2_ASAP7_75t_SL g640 ( 
.A(n_586),
.B(n_397),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_264),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_528),
.A2(n_422),
.B1(n_432),
.B2(n_426),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_559),
.B(n_463),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_526),
.B(n_459),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_525),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_572),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_538),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_582),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_569),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_525),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_525),
.B(n_465),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_551),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_554),
.B(n_447),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_551),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_582),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_553),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_556),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_556),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_539),
.B(n_512),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_576),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_579),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_560),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_547),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_531),
.B(n_343),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_R g676 ( 
.A(n_561),
.B(n_447),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_539),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_539),
.B(n_449),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_566),
.B(n_475),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_554),
.B(n_501),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_582),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_568),
.B(n_249),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_579),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_579),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_571),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_568),
.B(n_249),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_531),
.A2(n_292),
.B1(n_500),
.B2(n_460),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_541),
.B(n_345),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_586),
.B(n_211),
.Y(n_689)
);

CKINVDCx6p67_ASAP7_75t_R g690 ( 
.A(n_547),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_593),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_561),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_590),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_582),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_581),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_530),
.B(n_442),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_571),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_547),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_578),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_581),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_578),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_533),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_577),
.B(n_441),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_541),
.B(n_454),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_588),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_577),
.B(n_382),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_546),
.B(n_441),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_574),
.B(n_596),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_581),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_549),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_567),
.B(n_347),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_574),
.B(n_382),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_588),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_596),
.A2(n_323),
.B1(n_575),
.B2(n_567),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_580),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_549),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_549),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_549),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_517),
.Y(n_719)
);

AO22x1_ASAP7_75t_L g720 ( 
.A1(n_546),
.A2(n_230),
.B1(n_235),
.B2(n_229),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_575),
.B(n_382),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_583),
.B(n_461),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_588),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_562),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_590),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_535),
.B(n_263),
.C(n_262),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_549),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_535),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_R g732 ( 
.A(n_562),
.B(n_212),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_546),
.B(n_354),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_546),
.B(n_356),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_590),
.Y(n_735)
);

AO21x2_ASAP7_75t_L g736 ( 
.A1(n_550),
.A2(n_223),
.B(n_221),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_583),
.B(n_478),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_588),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_533),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_588),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_557),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_584),
.B(n_585),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_557),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_584),
.B(n_444),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_597),
.B(n_212),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_586),
.Y(n_747)
);

INVx11_ASAP7_75t_L g748 ( 
.A(n_540),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_537),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_557),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_715),
.B(n_587),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_691),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_743),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_743),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_612),
.B(n_264),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_646),
.A2(n_385),
.B1(n_260),
.B2(n_369),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_607),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_619),
.A2(n_247),
.B1(n_254),
.B2(n_226),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_640),
.B(n_264),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_640),
.B(n_267),
.Y(n_762)
);

AO221x1_ASAP7_75t_L g763 ( 
.A1(n_714),
.A2(n_337),
.B1(n_267),
.B2(n_265),
.C(n_257),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_715),
.B(n_726),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_726),
.B(n_587),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_SL g766 ( 
.A(n_728),
.B(n_230),
.C(n_229),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_608),
.B(n_216),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_750),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_708),
.B(n_587),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_640),
.A2(n_589),
.B1(n_267),
.B2(n_337),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_711),
.B(n_589),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_608),
.B(n_267),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_660),
.B(n_597),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_707),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_703),
.B(n_589),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_731),
.A2(n_589),
.B1(n_267),
.B2(n_337),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_604),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_679),
.B(n_216),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_607),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_647),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_707),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_645),
.B(n_337),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_644),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_521),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_645),
.B(n_521),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_645),
.B(n_337),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_737),
.A2(n_273),
.B1(n_335),
.B2(n_387),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_644),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_647),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_645),
.B(n_521),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_679),
.B(n_217),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_737),
.B(n_550),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_600),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_747),
.B(n_558),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_745),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_747),
.B(n_558),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_722),
.A2(n_359),
.B1(n_405),
.B2(n_242),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_644),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_660),
.B(n_496),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_675),
.B(n_273),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_745),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_604),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_599),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_656),
.B(n_599),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_648),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_605),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_738),
.A2(n_399),
.B1(n_238),
.B2(n_237),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_727),
.A2(n_735),
.B(n_693),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_704),
.B(n_466),
.C(n_458),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_680),
.B(n_217),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_656),
.B(n_565),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_610),
.B(n_565),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_610),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_615),
.B(n_537),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_601),
.B(n_658),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_688),
.A2(n_306),
.B1(n_274),
.B2(n_277),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_648),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_691),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_621),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_677),
.B(n_220),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_621),
.B(n_537),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_733),
.A2(n_542),
.B(n_533),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_693),
.B(n_273),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_642),
.B(n_220),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_600),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_687),
.A2(n_370),
.B1(n_325),
.B2(n_322),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_622),
.B(n_537),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_622),
.B(n_557),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_623),
.B(n_624),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_641),
.B(n_273),
.Y(n_832)
);

INVx4_ASAP7_75t_SL g833 ( 
.A(n_641),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_623),
.B(n_557),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_641),
.B(n_335),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_693),
.B(n_335),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_603),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_689),
.B(n_734),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_624),
.B(n_557),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_631),
.B(n_570),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_721),
.B(n_222),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_676),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_631),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_641),
.B(n_335),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_R g845 ( 
.A(n_732),
.B(n_552),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_649),
.B(n_496),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_222),
.Y(n_847)
);

BUFx5_ASAP7_75t_L g848 ( 
.A(n_727),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_632),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_692),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_639),
.A2(n_542),
.B(n_533),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_632),
.B(n_570),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_649),
.B(n_498),
.Y(n_853)
);

BUFx6f_ASAP7_75t_SL g854 ( 
.A(n_649),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_L g855 ( 
.A(n_641),
.B(n_335),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_686),
.B(n_227),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_706),
.A2(n_227),
.B1(n_232),
.B2(n_410),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_689),
.B(n_335),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_689),
.B(n_335),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_649),
.B(n_498),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_648),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_635),
.B(n_570),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_600),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_606),
.B(n_232),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_635),
.B(n_636),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_636),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_606),
.B(n_234),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_713),
.B(n_335),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_650),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_606),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_651),
.Y(n_871)
);

INVx4_ASAP7_75t_SL g872 ( 
.A(n_641),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_650),
.B(n_659),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_659),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_641),
.B(n_234),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_620),
.B(n_236),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_661),
.B(n_570),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_661),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_664),
.B(n_570),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_669),
.B(n_480),
.C(n_477),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_651),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_692),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_664),
.B(n_570),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_651),
.Y(n_884)
);

NOR2x1p5_ASAP7_75t_L g885 ( 
.A(n_690),
.B(n_235),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_634),
.B(n_236),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_665),
.B(n_237),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_665),
.B(n_545),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_667),
.B(n_545),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_667),
.B(n_536),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_674),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_696),
.B(n_392),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_668),
.B(n_672),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_678),
.B(n_238),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_602),
.B(n_241),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_725),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_613),
.B(n_585),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_713),
.B(n_279),
.Y(n_899)
);

NAND3xp33_ASAP7_75t_L g900 ( 
.A(n_609),
.B(n_746),
.C(n_712),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_672),
.A2(n_302),
.B1(n_283),
.B2(n_284),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_653),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_673),
.A2(n_390),
.B1(n_334),
.B2(n_317),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_617),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_673),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_685),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_685),
.B(n_536),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_SL g908 ( 
.A(n_735),
.B(n_533),
.Y(n_908)
);

OAI221xp5_ASAP7_75t_L g909 ( 
.A1(n_697),
.A2(n_482),
.B1(n_355),
.B2(n_373),
.C(n_300),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_748),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_697),
.B(n_536),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_699),
.A2(n_595),
.B1(n_594),
.B2(n_591),
.C(n_495),
.Y(n_912)
);

BUFx4_ASAP7_75t_L g913 ( 
.A(n_748),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_690),
.B(n_674),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_653),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_643),
.B(n_392),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_725),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_736),
.A2(n_595),
.B1(n_594),
.B2(n_591),
.Y(n_918)
);

OAI22x1_ASAP7_75t_SL g919 ( 
.A1(n_719),
.A2(n_376),
.B1(n_239),
.B2(n_383),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_699),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_713),
.B(n_241),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_617),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_764),
.B(n_701),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_808),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_757),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_753),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_817),
.B(n_701),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_842),
.B(n_638),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_817),
.B(n_638),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_776),
.A2(n_736),
.B1(n_392),
.B2(n_625),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_754),
.B(n_629),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_768),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_902),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_755),
.B(n_629),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_805),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_782),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_904),
.B(n_739),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_776),
.A2(n_638),
.B1(n_617),
.B2(n_749),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_813),
.B(n_736),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_815),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_915),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_814),
.B(n_749),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_795),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_752),
.B(n_749),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_821),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_795),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_774),
.A2(n_638),
.B1(n_628),
.B2(n_617),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_904),
.B(n_922),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_845),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_791),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_765),
.B(n_739),
.Y(n_951)
);

AND2x6_ASAP7_75t_L g952 ( 
.A(n_783),
.B(n_794),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_SL g953 ( 
.A(n_766),
.B(n_376),
.C(n_239),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_795),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_882),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_810),
.A2(n_455),
.B(n_495),
.C(n_493),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_843),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_849),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_775),
.B(n_739),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_866),
.Y(n_960)
);

INVx8_ASAP7_75t_L g961 ( 
.A(n_891),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_795),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_850),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_827),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_827),
.Y(n_965)
);

NOR2x1p5_ASAP7_75t_L g966 ( 
.A(n_910),
.B(n_383),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_827),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_827),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_820),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_895),
.A2(n_386),
.B1(n_393),
.B2(n_394),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_869),
.B(n_741),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_772),
.A2(n_618),
.B(n_684),
.C(n_695),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_874),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_878),
.B(n_741),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_896),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_905),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_797),
.B(n_616),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_906),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_922),
.B(n_741),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_767),
.B(n_720),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_L g981 ( 
.A(n_770),
.B(n_702),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_SL g982 ( 
.A1(n_897),
.A2(n_386),
.B1(n_393),
.B2(n_394),
.Y(n_982)
);

AND2x4_ASAP7_75t_SL g983 ( 
.A(n_777),
.B(n_674),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_804),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_863),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_770),
.A2(n_694),
.B1(n_681),
.B2(n_705),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_778),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_863),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_803),
.B(n_773),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_761),
.A2(n_611),
.B1(n_614),
.B2(n_700),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_917),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_898),
.B(n_451),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_863),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_920),
.B(n_603),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_890),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_831),
.B(n_603),
.Y(n_996)
);

AND2x6_ASAP7_75t_SL g997 ( 
.A(n_895),
.B(n_455),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_845),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_863),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_846),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_907),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_780),
.A2(n_467),
.B(n_493),
.C(n_491),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_853),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_900),
.A2(n_694),
.B1(n_681),
.B2(n_705),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_865),
.B(n_603),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_778),
.B(n_654),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_759),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_860),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_870),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_838),
.A2(n_740),
.B(n_702),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_870),
.B(n_654),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_911),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_848),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_806),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_848),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_891),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_801),
.B(n_457),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_767),
.B(n_720),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_916),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_816),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_848),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_873),
.B(n_654),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_779),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_771),
.A2(n_694),
.B1(n_681),
.B2(n_705),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_893),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_823),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_761),
.A2(n_627),
.B1(n_630),
.B2(n_611),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_892),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_829),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_830),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_SL g1031 ( 
.A1(n_908),
.A2(n_723),
.B(n_705),
.C(n_681),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_848),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_780),
.B(n_654),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_793),
.B(n_694),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_834),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_913),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_822),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_769),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_793),
.B(n_772),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_826),
.B(n_723),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_839),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_781),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_848),
.B(n_674),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_785),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_762),
.A2(n_630),
.B1(n_633),
.B2(n_614),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_840),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_786),
.A2(n_723),
.B1(n_729),
.B2(n_724),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_888),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_852),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_854),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_812),
.B(n_723),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_833),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_SL g1053 ( 
.A1(n_762),
.A2(n_467),
.B(n_457),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_796),
.B(n_729),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_880),
.B(n_468),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_862),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_790),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_800),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_812),
.B(n_729),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_841),
.A2(n_729),
.B1(n_751),
.B2(n_724),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_877),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_879),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_833),
.B(n_468),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_883),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_798),
.A2(n_398),
.B1(n_409),
.B2(n_326),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_825),
.A2(n_716),
.B(n_710),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_889),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_807),
.B(n_742),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_914),
.B(n_698),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_848),
.B(n_698),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_819),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_809),
.B(n_822),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_864),
.B(n_710),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_919),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_861),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_838),
.B(n_698),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_871),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_841),
.A2(n_751),
.B1(n_716),
.B2(n_717),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_884),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_868),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_868),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_864),
.B(n_867),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_837),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_867),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_825),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_899),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_836),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_876),
.A2(n_698),
.B1(n_398),
.B2(n_379),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_787),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_918),
.B(n_717),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_899),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_912),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_847),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_789),
.A2(n_618),
.B1(n_625),
.B2(n_626),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_836),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_833),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_854),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_802),
.A2(n_718),
.B(n_730),
.C(n_744),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_847),
.A2(n_718),
.B1(n_730),
.B2(n_744),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_918),
.B(n_742),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_SL g1103 ( 
.A(n_828),
.B(n_269),
.C(n_266),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_872),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_789),
.B(n_742),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_921),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_792),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_894),
.B(n_744),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_856),
.A2(n_242),
.B1(n_400),
.B2(n_374),
.Y(n_1109)
);

AO22x1_ASAP7_75t_L g1110 ( 
.A1(n_876),
.A2(n_311),
.B1(n_297),
.B2(n_295),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_856),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_802),
.Y(n_1112)
);

AND3x2_ASAP7_75t_SL g1113 ( 
.A(n_886),
.B(n_0),
.C(n_1),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_872),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_799),
.B(n_278),
.C(n_270),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_926),
.B(n_894),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_943),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_923),
.B(n_886),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_981),
.A2(n_788),
.B(n_784),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_925),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1072),
.A2(n_1037),
.B1(n_980),
.B2(n_1018),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_961),
.B(n_921),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_925),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1072),
.A2(n_818),
.B1(n_760),
.B2(n_763),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_SL g1125 ( 
.A(n_929),
.B(n_909),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1094),
.B(n_758),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_948),
.A2(n_788),
.B(n_784),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_932),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_948),
.A2(n_859),
.B(n_858),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1076),
.A2(n_859),
.B(n_858),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_943),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_932),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_955),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_923),
.B(n_811),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_927),
.B(n_887),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1019),
.A2(n_857),
.B1(n_341),
.B2(n_371),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_987),
.A2(n_756),
.B(n_824),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_945),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_929),
.B(n_1052),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1083),
.B(n_756),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_989),
.B(n_872),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_987),
.A2(n_875),
.B(n_835),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_989),
.B(n_469),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1028),
.B(n_901),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1077),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1039),
.A2(n_855),
.B(n_844),
.C(n_832),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_949),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_943),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_945),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1028),
.B(n_903),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_987),
.A2(n_662),
.B(n_652),
.Y(n_1151)
);

BUFx4f_ASAP7_75t_L g1152 ( 
.A(n_961),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_987),
.A2(n_938),
.B(n_1015),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1085),
.A2(n_374),
.B1(n_410),
.B2(n_379),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_1016),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1094),
.B(n_389),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1102),
.A2(n_851),
.B(n_709),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1054),
.A2(n_652),
.B(n_662),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_951),
.A2(n_652),
.B(n_662),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1115),
.B(n_308),
.C(n_286),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_944),
.A2(n_652),
.B(n_662),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1065),
.A2(n_474),
.B(n_470),
.C(n_472),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1065),
.A2(n_474),
.B(n_470),
.C(n_472),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_943),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_930),
.A2(n_301),
.B1(n_315),
.B2(n_319),
.Y(n_1165)
);

O2A1O1Ixp5_ASAP7_75t_L g1166 ( 
.A1(n_1076),
.A2(n_627),
.B(n_626),
.C(n_633),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_959),
.A2(n_652),
.B(n_662),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_962),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_962),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_973),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_962),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1002),
.A2(n_469),
.B(n_483),
.C(n_484),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_982),
.B(n_333),
.C(n_329),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_998),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1102),
.A2(n_637),
.B(n_684),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1111),
.B(n_321),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1111),
.B(n_389),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1000),
.B(n_1003),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_955),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1000),
.B(n_395),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1050),
.B(n_324),
.C(n_336),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1110),
.B(n_346),
.C(n_365),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1079),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1105),
.A2(n_652),
.B(n_662),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1003),
.B(n_395),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_962),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1106),
.A2(n_400),
.B(n_399),
.C(n_396),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1009),
.A2(n_740),
.B(n_702),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1008),
.B(n_483),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1025),
.B(n_637),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1008),
.B(n_931),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1025),
.A2(n_396),
.B(n_695),
.C(n_700),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1073),
.A2(n_653),
.B(n_709),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1079),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1016),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_924),
.B(n_702),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_936),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_930),
.A2(n_338),
.B1(n_342),
.B2(n_350),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1014),
.B(n_655),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1051),
.A2(n_353),
.B(n_401),
.C(n_357),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_973),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_936),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1109),
.A2(n_358),
.B1(n_363),
.B2(n_360),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_926),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1051),
.A2(n_361),
.B(n_403),
.C(n_709),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1080),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1014),
.B(n_655),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_984),
.B(n_702),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1002),
.A2(n_491),
.B(n_484),
.C(n_487),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1059),
.A2(n_657),
.B(n_655),
.C(n_683),
.Y(n_1210)
);

OAI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1074),
.A2(n_487),
.B1(n_488),
.B2(n_490),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_963),
.B(n_991),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1048),
.B(n_702),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1048),
.A2(n_490),
.B(n_488),
.C(n_657),
.Y(n_1214)
);

AOI22x1_ASAP7_75t_L g1215 ( 
.A1(n_995),
.A2(n_657),
.B1(n_683),
.B2(n_671),
.Y(n_1215)
);

OR2x6_ASAP7_75t_SL g1216 ( 
.A(n_1099),
.B(n_444),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_975),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1052),
.B(n_663),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_975),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1067),
.B(n_663),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_931),
.B(n_68),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1080),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1009),
.A2(n_740),
.B(n_533),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1067),
.B(n_663),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_969),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1059),
.A2(n_666),
.B(n_683),
.C(n_671),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1089),
.B(n_494),
.C(n_514),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1040),
.A2(n_671),
.B(n_670),
.C(n_666),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_928),
.A2(n_740),
.B1(n_670),
.B2(n_666),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_984),
.B(n_740),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1001),
.B(n_670),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_934),
.B(n_137),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_935),
.Y(n_1233)
);

AO32x1_ASAP7_75t_L g1234 ( 
.A1(n_986),
.A2(n_514),
.A3(n_494),
.B1(n_7),
.B2(n_11),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1093),
.A2(n_956),
.B(n_1053),
.C(n_928),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_940),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_950),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1091),
.A2(n_740),
.B1(n_5),
.B2(n_15),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1017),
.B(n_0),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_956),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1012),
.B(n_16),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1030),
.B(n_542),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_942),
.A2(n_542),
.B(n_206),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1086),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_996),
.A2(n_542),
.B(n_79),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1086),
.A2(n_1088),
.B1(n_1096),
.B2(n_978),
.Y(n_1246)
);

O2A1O1Ixp5_ASAP7_75t_SL g1247 ( 
.A1(n_1108),
.A2(n_958),
.B(n_960),
.C(n_957),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_969),
.B(n_21),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_976),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1103),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_933),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_933),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_941),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1017),
.B(n_22),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1035),
.B(n_27),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1041),
.B(n_28),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_941),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1075),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_971),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1055),
.A2(n_31),
.B(n_34),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1088),
.A2(n_1096),
.B1(n_1032),
.B2(n_1013),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1005),
.A2(n_542),
.B(n_104),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_977),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1022),
.A2(n_98),
.B(n_195),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1046),
.B(n_38),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_937),
.A2(n_94),
.B(n_188),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1040),
.A2(n_38),
.B(n_39),
.C(n_41),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_R g1268 ( 
.A(n_961),
.B(n_106),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1103),
.A2(n_43),
.B(n_47),
.C(n_48),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1013),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_997),
.B(n_52),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_992),
.B(n_53),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_974),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1049),
.B(n_54),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_947),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_993),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1038),
.A2(n_55),
.B(n_60),
.C(n_64),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_937),
.A2(n_979),
.B(n_1021),
.Y(n_1278)
);

CKINVDCx12_ASAP7_75t_R g1279 ( 
.A(n_1122),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1118),
.B(n_1056),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1168),
.B(n_999),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1119),
.A2(n_1043),
.B(n_1070),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1233),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1137),
.A2(n_1043),
.B(n_1070),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1132),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1175),
.A2(n_1010),
.B(n_1100),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1278),
.A2(n_1066),
.B(n_972),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1235),
.A2(n_1021),
.B(n_1032),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1210),
.A2(n_939),
.B(n_1033),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1157),
.A2(n_1006),
.B(n_979),
.Y(n_1290)
);

NAND2x1_ASAP7_75t_L g1291 ( 
.A(n_1168),
.B(n_964),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1129),
.A2(n_1034),
.B(n_1090),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_953),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1153),
.A2(n_1090),
.B(n_1107),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1238),
.A2(n_1064),
.B1(n_1062),
.B2(n_1061),
.C(n_1026),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1126),
.A2(n_1055),
.B(n_1113),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1237),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1157),
.A2(n_1006),
.B(n_994),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1143),
.B(n_953),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1134),
.B(n_1038),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1236),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1259),
.B(n_992),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1193),
.A2(n_1004),
.B(n_1011),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1273),
.B(n_1020),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1204),
.Y(n_1305)
);

NAND2x1_ASAP7_75t_L g1306 ( 
.A(n_1186),
.B(n_964),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1127),
.A2(n_1218),
.B(n_1146),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1145),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1130),
.A2(n_1011),
.B(n_1112),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1189),
.B(n_977),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1166),
.A2(n_1045),
.B(n_1027),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1260),
.A2(n_934),
.B1(n_952),
.B2(n_1087),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1226),
.A2(n_1078),
.B(n_1101),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1147),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1225),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1135),
.B(n_1029),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1215),
.A2(n_1027),
.B(n_990),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1140),
.A2(n_993),
.B(n_1090),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1142),
.A2(n_1107),
.B(n_954),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1152),
.B(n_1036),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1165),
.A2(n_970),
.B1(n_1098),
.B2(n_1036),
.C(n_1092),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1121),
.A2(n_952),
.B1(n_966),
.B2(n_1063),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1125),
.A2(n_952),
.B1(n_1082),
.B2(n_1063),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1133),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1212),
.B(n_983),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1125),
.A2(n_1060),
.B(n_1081),
.C(n_983),
.Y(n_1326)
);

AO32x2_ASAP7_75t_L g1327 ( 
.A1(n_1238),
.A2(n_1113),
.A3(n_985),
.B1(n_968),
.B2(n_952),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1131),
.Y(n_1328)
);

AOI211x1_ASAP7_75t_L g1329 ( 
.A1(n_1275),
.A2(n_1084),
.B(n_952),
.C(n_65),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1176),
.B(n_1116),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1124),
.B(n_1024),
.C(n_1047),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1189),
.B(n_1007),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1225),
.B(n_1069),
.Y(n_1333)
);

AOI21xp33_ASAP7_75t_L g1334 ( 
.A1(n_1250),
.A2(n_1107),
.B(n_1031),
.Y(n_1334)
);

OA22x2_ASAP7_75t_L g1335 ( 
.A1(n_1211),
.A2(n_1081),
.B1(n_1104),
.B2(n_1097),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1249),
.B(n_999),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1184),
.A2(n_990),
.B(n_1045),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1228),
.A2(n_1095),
.B(n_1031),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1261),
.A2(n_968),
.B(n_985),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1261),
.A2(n_1095),
.B(n_946),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1267),
.A2(n_1023),
.B(n_1058),
.C(n_1057),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1178),
.B(n_946),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_1248),
.Y(n_1343)
);

AO21x1_ASAP7_75t_L g1344 ( 
.A1(n_1269),
.A2(n_1114),
.B(n_1104),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_SL g1345 ( 
.A1(n_1205),
.A2(n_1114),
.B(n_1097),
.C(n_965),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1139),
.A2(n_993),
.B(n_1071),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1241),
.B(n_965),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1199),
.B(n_967),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1152),
.B(n_993),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1161),
.A2(n_967),
.B(n_988),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1246),
.A2(n_1042),
.B(n_1069),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1239),
.B(n_988),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1158),
.A2(n_1058),
.B(n_1057),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1139),
.A2(n_1071),
.B(n_1042),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_SL g1355 ( 
.A1(n_1255),
.A2(n_1068),
.B(n_1071),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1120),
.A2(n_1071),
.B1(n_1044),
.B2(n_1023),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1188),
.A2(n_1042),
.B(n_1044),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1223),
.A2(n_1068),
.B(n_1042),
.Y(n_1358)
);

O2A1O1Ixp5_ASAP7_75t_L g1359 ( 
.A1(n_1144),
.A2(n_1068),
.B(n_91),
.C(n_115),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1131),
.Y(n_1360)
);

AO32x2_ASAP7_75t_L g1361 ( 
.A1(n_1244),
.A2(n_1068),
.A3(n_118),
.B1(n_120),
.B2(n_126),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1179),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1207),
.B(n_1220),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1174),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1123),
.A2(n_1217),
.B1(n_1149),
.B2(n_1201),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1224),
.B(n_1068),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1128),
.B(n_81),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1159),
.A2(n_130),
.B(n_140),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1138),
.B(n_143),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1246),
.A2(n_148),
.B(n_158),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1245),
.A2(n_164),
.B(n_177),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1141),
.B(n_185),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1197),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1141),
.B(n_186),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1170),
.B(n_198),
.Y(n_1375)
);

OAI22x1_ASAP7_75t_L g1376 ( 
.A1(n_1271),
.A2(n_1150),
.B1(n_1177),
.B2(n_1156),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1219),
.B(n_1190),
.Y(n_1377)
);

INVx3_ASAP7_75t_SL g1378 ( 
.A(n_1202),
.Y(n_1378)
);

AOI221x1_ASAP7_75t_L g1379 ( 
.A1(n_1244),
.A2(n_1270),
.B1(n_1243),
.B2(n_1262),
.C(n_1277),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1200),
.A2(n_1160),
.B(n_1274),
.C(n_1265),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1263),
.B(n_1191),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1231),
.A2(n_1167),
.B(n_1242),
.Y(n_1382)
);

CKINVDCx6p67_ASAP7_75t_R g1383 ( 
.A(n_1195),
.Y(n_1383)
);

BUFx10_ASAP7_75t_L g1384 ( 
.A(n_1272),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1203),
.B(n_1185),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1256),
.A2(n_1192),
.B(n_1240),
.C(n_1227),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1247),
.A2(n_1242),
.B(n_1151),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1258),
.B(n_1213),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1270),
.A2(n_1187),
.A3(n_1264),
.B(n_1257),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1208),
.A2(n_1230),
.B(n_1164),
.Y(n_1390)
);

NOR2x1_ASAP7_75t_L g1391 ( 
.A(n_1186),
.B(n_1117),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1229),
.A2(n_1266),
.B(n_1253),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1196),
.A2(n_1234),
.B(n_1180),
.Y(n_1393)
);

OAI21xp33_ASAP7_75t_L g1394 ( 
.A1(n_1165),
.A2(n_1198),
.B(n_1154),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1131),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1191),
.B(n_1254),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1183),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1194),
.Y(n_1398)
);

OAI22x1_ASAP7_75t_L g1399 ( 
.A1(n_1221),
.A2(n_1232),
.B1(n_1222),
.B2(n_1206),
.Y(n_1399)
);

AO21x1_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1182),
.B(n_1198),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1221),
.A2(n_1232),
.B1(n_1136),
.B2(n_1122),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1122),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1209),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1148),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1234),
.A2(n_1173),
.B(n_1181),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1117),
.B(n_1169),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1268),
.B(n_1148),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1172),
.A2(n_1169),
.B(n_1234),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1148),
.A2(n_1171),
.B(n_1276),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1171),
.A2(n_1276),
.B(n_1216),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1171),
.A2(n_1276),
.B(n_1072),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1118),
.B(n_1134),
.Y(n_1413)
);

AO21x1_ASAP7_75t_L g1414 ( 
.A1(n_1118),
.A2(n_1238),
.B(n_1083),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1118),
.B(n_1134),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1417)
);

AO32x2_ASAP7_75t_L g1418 ( 
.A1(n_1238),
.A2(n_1244),
.A3(n_1270),
.B1(n_1261),
.B2(n_1246),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1118),
.A2(n_776),
.B1(n_764),
.B2(n_770),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1153),
.A2(n_1076),
.B(n_1193),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1118),
.B(n_923),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1212),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1233),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1212),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1216),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1141),
.B(n_1191),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1153),
.A2(n_1076),
.B(n_1193),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1175),
.A2(n_1278),
.B(n_1010),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1155),
.Y(n_1430)
);

AO32x2_ASAP7_75t_L g1431 ( 
.A1(n_1238),
.A2(n_1244),
.A3(n_1270),
.B1(n_1261),
.B2(n_1246),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1175),
.A2(n_1278),
.B(n_1010),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1132),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1134),
.B(n_1028),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1143),
.B(n_980),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1233),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_SL g1439 ( 
.A(n_1152),
.B(n_854),
.Y(n_1439)
);

NAND3x1_ASAP7_75t_L g1440 ( 
.A(n_1271),
.B(n_1113),
.C(n_696),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1118),
.B(n_1134),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1233),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1118),
.A2(n_776),
.B1(n_764),
.B2(n_770),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1131),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1118),
.A2(n_776),
.B1(n_764),
.B2(n_770),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1204),
.Y(n_1446)
);

AO31x2_ASAP7_75t_L g1447 ( 
.A1(n_1121),
.A2(n_1261),
.A3(n_1226),
.B(n_1119),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1132),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1119),
.A2(n_922),
.B(n_904),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1437),
.B(n_1330),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_SL g1452 ( 
.A1(n_1380),
.A2(n_1386),
.B(n_1394),
.C(n_1445),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1295),
.A2(n_1387),
.B(n_1379),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1307),
.A2(n_1428),
.B(n_1420),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1284),
.A2(n_1289),
.B(n_1282),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1456)
);

OAI222xp33_ASAP7_75t_L g1457 ( 
.A1(n_1312),
.A2(n_1415),
.B1(n_1413),
.B2(n_1441),
.C1(n_1401),
.C2(n_1300),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1382),
.A2(n_1303),
.B(n_1292),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1350),
.A2(n_1417),
.B(n_1416),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1424),
.A2(n_1433),
.B(n_1432),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1308),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1421),
.B(n_1280),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1394),
.A2(n_1385),
.B1(n_1414),
.B2(n_1421),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1310),
.B(n_1332),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1400),
.A2(n_1404),
.B1(n_1376),
.B2(n_1436),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1449),
.A2(n_1309),
.B(n_1353),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1351),
.B(n_1318),
.Y(n_1467)
);

AOI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1404),
.A2(n_1443),
.B(n_1419),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1397),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1419),
.A2(n_1443),
.B1(n_1445),
.B2(n_1331),
.Y(n_1470)
);

NOR2xp67_ASAP7_75t_L g1471 ( 
.A(n_1425),
.B(n_1314),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1422),
.B(n_1396),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1305),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1285),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1315),
.B(n_1297),
.Y(n_1476)
);

AND2x6_ASAP7_75t_L g1477 ( 
.A(n_1323),
.B(n_1312),
.Y(n_1477)
);

INVxp33_ASAP7_75t_L g1478 ( 
.A(n_1381),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1293),
.B(n_1299),
.Y(n_1479)
);

AO221x2_ASAP7_75t_L g1480 ( 
.A1(n_1296),
.A2(n_1440),
.B1(n_1409),
.B2(n_1361),
.C(n_1327),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1287),
.A2(n_1290),
.B(n_1337),
.Y(n_1481)
);

AOI31xp67_ASAP7_75t_L g1482 ( 
.A1(n_1323),
.A2(n_1335),
.A3(n_1401),
.B(n_1366),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1483)
);

NOR2xp67_ASAP7_75t_L g1484 ( 
.A(n_1364),
.B(n_1325),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1405),
.B(n_1315),
.Y(n_1485)
);

AOI221x1_ASAP7_75t_L g1486 ( 
.A1(n_1334),
.A2(n_1393),
.B1(n_1370),
.B2(n_1409),
.C(n_1412),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1283),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1304),
.B(n_1316),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1368),
.A2(n_1355),
.B(n_1298),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1392),
.A2(n_1294),
.B(n_1358),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1331),
.A2(n_1321),
.B1(n_1343),
.B2(n_1406),
.Y(n_1491)
);

NAND2x1_ASAP7_75t_L g1492 ( 
.A(n_1288),
.B(n_1354),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1352),
.B(n_1427),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1319),
.A2(n_1317),
.B(n_1340),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1295),
.A2(n_1289),
.B(n_1334),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1373),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1447),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1344),
.A2(n_1346),
.B(n_1341),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1435),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1296),
.A2(n_1326),
.B(n_1302),
.C(n_1359),
.Y(n_1500)
);

AOI21xp33_ASAP7_75t_L g1501 ( 
.A1(n_1347),
.A2(n_1399),
.B(n_1388),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1311),
.A2(n_1339),
.B(n_1357),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1448),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1378),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1301),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1371),
.A2(n_1365),
.B(n_1338),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1338),
.A2(n_1313),
.B(n_1356),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1345),
.A2(n_1363),
.B(n_1377),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1423),
.B(n_1438),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1442),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1430),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1313),
.A2(n_1356),
.B(n_1390),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1427),
.B(n_1398),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1402),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1377),
.B(n_1342),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1412),
.A2(n_1348),
.B(n_1375),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1324),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1405),
.B(n_1403),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1410),
.A2(n_1369),
.B(n_1367),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1322),
.A2(n_1407),
.B(n_1291),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1306),
.A2(n_1391),
.B(n_1336),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1395),
.Y(n_1522)
);

AOI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1333),
.A2(n_1406),
.B(n_1408),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1447),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1281),
.A2(n_1395),
.B(n_1411),
.Y(n_1525)
);

AO31x2_ASAP7_75t_L g1526 ( 
.A1(n_1418),
.A2(n_1431),
.A3(n_1327),
.B(n_1447),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1281),
.A2(n_1320),
.B(n_1349),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1389),
.A2(n_1418),
.B(n_1431),
.Y(n_1528)
);

AOI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1418),
.A2(n_1431),
.B(n_1389),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1343),
.B(n_1384),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1361),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1361),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1328),
.B(n_1444),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1349),
.A2(n_1320),
.B(n_1439),
.C(n_1327),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1328),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1329),
.B(n_1362),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1384),
.B(n_1439),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1444),
.Y(n_1538)
);

O2A1O1Ixp5_ASAP7_75t_L g1539 ( 
.A1(n_1279),
.A2(n_1405),
.B(n_1360),
.C(n_1444),
.Y(n_1539)
);

BUFx2_ASAP7_75t_SL g1540 ( 
.A(n_1360),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1383),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1426),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1330),
.A2(n_1118),
.B1(n_1028),
.B2(n_1072),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1372),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1351),
.B(n_1318),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1394),
.A2(n_1118),
.B1(n_1072),
.B2(n_1134),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1372),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1314),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1373),
.Y(n_1554)
);

AOI22x1_ASAP7_75t_L g1555 ( 
.A1(n_1376),
.A2(n_1085),
.B1(n_1121),
.B2(n_1399),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1385),
.A2(n_1072),
.B1(n_1394),
.B2(n_413),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1416),
.A2(n_981),
.B(n_1417),
.Y(n_1557)
);

XNOR2xp5_ASAP7_75t_L g1558 ( 
.A(n_1364),
.B(n_517),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1373),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1308),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1308),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_1414),
.A2(n_1118),
.B(n_1344),
.C(n_1028),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1394),
.A2(n_1118),
.B(n_1072),
.C(n_1134),
.Y(n_1569)
);

BUFx2_ASAP7_75t_R g1570 ( 
.A(n_1314),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_SL g1572 ( 
.A1(n_1380),
.A2(n_1267),
.B(n_1118),
.C(n_1386),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1308),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1394),
.A2(n_1118),
.B(n_1072),
.C(n_1134),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1373),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1295),
.A2(n_1387),
.B(n_1379),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1283),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1446),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1394),
.A2(n_1118),
.B(n_1072),
.C(n_1419),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1394),
.A2(n_1118),
.B(n_1072),
.C(n_1419),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1420),
.A2(n_1193),
.B(n_1428),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1330),
.A2(n_949),
.B(n_1271),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1283),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1394),
.A2(n_1118),
.B1(n_1072),
.B2(n_1134),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1592)
);

AO21x1_ASAP7_75t_L g1593 ( 
.A1(n_1296),
.A2(n_1238),
.B(n_1118),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1283),
.Y(n_1594)
);

INVx3_ASAP7_75t_SL g1595 ( 
.A(n_1314),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_SL g1597 ( 
.A1(n_1400),
.A2(n_1344),
.B(n_1404),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1598)
);

AOI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1420),
.A2(n_1193),
.B(n_1428),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1283),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1283),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1437),
.B(n_1330),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1295),
.A2(n_1387),
.B(n_1379),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1308),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1308),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1437),
.B(n_1330),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1608)
);

AOI22x1_ASAP7_75t_L g1609 ( 
.A1(n_1376),
.A2(n_1085),
.B1(n_1121),
.B2(n_1399),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1413),
.A2(n_1118),
.B(n_1072),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1296),
.A2(n_1118),
.B1(n_1134),
.B2(n_1413),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1283),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1286),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1485),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1486),
.A2(n_1454),
.B(n_1507),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1545),
.B(n_1567),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1487),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1545),
.B(n_1567),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1474),
.B(n_1478),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1524),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1454),
.A2(n_1507),
.B(n_1506),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1451),
.B(n_1602),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1556),
.A2(n_1549),
.B1(n_1591),
.B2(n_1571),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1607),
.B(n_1479),
.Y(n_1627)
);

NOR2xp67_ASAP7_75t_L g1628 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1628)
);

NOR2xp67_ASAP7_75t_L g1629 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1569),
.A2(n_1575),
.B(n_1580),
.C(n_1582),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1473),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1549),
.A2(n_1591),
.B1(n_1590),
.B2(n_1571),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1580),
.A2(n_1582),
.B(n_1572),
.C(n_1543),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1505),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1583),
.A2(n_1590),
.B1(n_1598),
.B2(n_1547),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1478),
.B(n_1464),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1494),
.A2(n_1502),
.B(n_1468),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1572),
.A2(n_1612),
.B(n_1611),
.C(n_1452),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1493),
.B(n_1513),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1513),
.B(n_1583),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1463),
.B(n_1465),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1546),
.B(n_1488),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1456),
.B(n_1483),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1456),
.B(n_1483),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1463),
.A2(n_1534),
.B(n_1465),
.C(n_1566),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1504),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1510),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1485),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1578),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1462),
.A2(n_1491),
.B1(n_1610),
.B2(n_1613),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1579),
.Y(n_1651)
);

AOI21x1_ASAP7_75t_SL g1652 ( 
.A1(n_1537),
.A2(n_1515),
.B(n_1533),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1595),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1514),
.B(n_1461),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1586),
.B(n_1610),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1496),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1570),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1588),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1586),
.B(n_1610),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1595),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1594),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1467),
.A2(n_1548),
.B(n_1452),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1600),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1601),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1461),
.B(n_1469),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1491),
.A2(n_1613),
.B1(n_1551),
.B2(n_1544),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1509),
.B(n_1614),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1469),
.B(n_1475),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1480),
.B(n_1475),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1467),
.A2(n_1548),
.B(n_1508),
.Y(n_1670)
);

O2A1O1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1457),
.A2(n_1500),
.B(n_1585),
.C(n_1597),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1544),
.B(n_1551),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1536),
.A2(n_1500),
.B1(n_1470),
.B2(n_1484),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1533),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1536),
.A2(n_1470),
.B1(n_1471),
.B2(n_1548),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1467),
.A2(n_1557),
.B(n_1455),
.Y(n_1677)
);

O2A1O1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1593),
.A2(n_1501),
.B(n_1498),
.C(n_1527),
.Y(n_1678)
);

AOI21x1_ASAP7_75t_SL g1679 ( 
.A1(n_1480),
.A2(n_1555),
.B(n_1609),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1562),
.B(n_1565),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1534),
.A2(n_1516),
.B(n_1558),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1492),
.A2(n_1495),
.B(n_1458),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1517),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1565),
.B(n_1574),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1604),
.B(n_1605),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1477),
.B(n_1522),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1518),
.A2(n_1504),
.B1(n_1576),
.B2(n_1554),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1518),
.A2(n_1561),
.B1(n_1541),
.B2(n_1523),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1477),
.B(n_1538),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1512),
.A2(n_1458),
.B(n_1481),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1477),
.B(n_1516),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1511),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1516),
.B(n_1526),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1535),
.B(n_1540),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1482),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1696)
);

AOI21x1_ASAP7_75t_SL g1697 ( 
.A1(n_1453),
.A2(n_1603),
.B(n_1577),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1477),
.B(n_1526),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1477),
.B(n_1526),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1525),
.B(n_1521),
.Y(n_1700)
);

OR2x6_ASAP7_75t_L g1701 ( 
.A(n_1512),
.B(n_1520),
.Y(n_1701)
);

CKINVDCx16_ASAP7_75t_R g1702 ( 
.A(n_1511),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1495),
.A2(n_1460),
.B(n_1459),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1497),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1521),
.B(n_1520),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1495),
.A2(n_1460),
.B(n_1459),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1707)
);

O2A1O1Ixp5_ASAP7_75t_L g1708 ( 
.A1(n_1529),
.A2(n_1584),
.B(n_1599),
.C(n_1532),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1481),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1542),
.A2(n_1531),
.B1(n_1453),
.B2(n_1577),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1489),
.B(n_1519),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1577),
.B(n_1603),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1531),
.B(n_1603),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1542),
.B(n_1519),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1542),
.B(n_1490),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1490),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1450),
.A2(n_1573),
.B(n_1550),
.C(n_1552),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1559),
.A2(n_1587),
.B(n_1560),
.C(n_1563),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1466),
.A2(n_1563),
.B1(n_1564),
.B2(n_1568),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1581),
.A2(n_1587),
.B(n_1589),
.C(n_1592),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1589),
.A2(n_1592),
.B(n_1596),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1596),
.A2(n_1606),
.B(n_1608),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1615),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1615),
.B(n_1545),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1486),
.A2(n_1295),
.B(n_1454),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1487),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1569),
.A2(n_1118),
.B(n_981),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1556),
.A2(n_1591),
.B1(n_1549),
.B2(n_1394),
.C(n_1028),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1451),
.B(n_1602),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1556),
.A2(n_1440),
.B1(n_1591),
.B2(n_1549),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1556),
.A2(n_1440),
.B1(n_1591),
.B2(n_1549),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1545),
.B(n_1567),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1569),
.A2(n_1575),
.B(n_1582),
.C(n_1580),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1485),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1487),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1486),
.A2(n_1295),
.B(n_1454),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1487),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1740)
);

NOR2xp67_ASAP7_75t_L g1741 ( 
.A(n_1553),
.B(n_1016),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1487),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1569),
.A2(n_1575),
.B(n_1118),
.C(n_1556),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1451),
.B(n_1602),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1451),
.B(n_1602),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1703),
.A2(n_1706),
.B(n_1682),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1707),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1693),
.B(n_1714),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1623),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1705),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1711),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1698),
.B(n_1699),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1691),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1677),
.A2(n_1720),
.B(n_1719),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1634),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1726),
.B(n_1669),
.Y(n_1758)
);

OR2x6_ASAP7_75t_L g1759 ( 
.A(n_1670),
.B(n_1701),
.Y(n_1759)
);

BUFx4f_ASAP7_75t_SL g1760 ( 
.A(n_1660),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1708),
.A2(n_1720),
.B(n_1719),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1704),
.B(n_1727),
.Y(n_1762)
);

BUFx4f_ASAP7_75t_SL g1763 ( 
.A(n_1660),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1697),
.A2(n_1722),
.B(n_1721),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1712),
.Y(n_1766)
);

AO21x2_ASAP7_75t_L g1767 ( 
.A1(n_1724),
.A2(n_1696),
.B(n_1718),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1732),
.A2(n_1733),
.B1(n_1730),
.B2(n_1641),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1710),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1647),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1701),
.B(n_1717),
.Y(n_1771)
);

AOI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1641),
.A2(n_1662),
.B(n_1688),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_R g1773 ( 
.A(n_1657),
.B(n_1692),
.Y(n_1773)
);

OA21x2_ASAP7_75t_L g1774 ( 
.A1(n_1645),
.A2(n_1725),
.B(n_1695),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1618),
.B(n_1738),
.Y(n_1775)
);

CKINVDCx11_ASAP7_75t_R g1776 ( 
.A(n_1702),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1621),
.B(n_1734),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1658),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1642),
.B(n_1658),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1716),
.B(n_1715),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1620),
.Y(n_1781)
);

OAI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1743),
.A2(n_1735),
.B(n_1630),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1723),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1715),
.B(n_1637),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1686),
.A2(n_1743),
.B(n_1729),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1689),
.A2(n_1728),
.B(n_1649),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1661),
.Y(n_1787)
);

AO21x2_ASAP7_75t_L g1788 ( 
.A1(n_1681),
.A2(n_1678),
.B(n_1673),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1663),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1633),
.A2(n_1650),
.B(n_1666),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1664),
.B(n_1737),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1739),
.B(n_1742),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1680),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1665),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1616),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1668),
.Y(n_1797)
);

AO21x2_ASAP7_75t_L g1798 ( 
.A1(n_1697),
.A2(n_1676),
.B(n_1671),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1624),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1674),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1636),
.A2(n_1622),
.B1(n_1627),
.B2(n_1744),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1684),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1616),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1755),
.B(n_1617),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1771),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1747),
.B(n_1690),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1764),
.B(n_1656),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1778),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1747),
.B(n_1640),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1771),
.Y(n_1810)
);

NOR2x1p5_ASAP7_75t_L g1811 ( 
.A(n_1772),
.B(n_1648),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1784),
.B(n_1685),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1755),
.B(n_1800),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1800),
.B(n_1740),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1752),
.B(n_1745),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1757),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1748),
.B(n_1667),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1783),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1752),
.B(n_1625),
.Y(n_1819)
);

NAND2x1p5_ASAP7_75t_L g1820 ( 
.A(n_1761),
.B(n_1648),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1748),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1764),
.A2(n_1638),
.B1(n_1683),
.B2(n_1631),
.C(n_1651),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1748),
.B(n_1654),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1753),
.B(n_1736),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1783),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1786),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1769),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1753),
.B(n_1736),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1746),
.A2(n_1679),
.B(n_1652),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1753),
.B(n_1731),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1751),
.B(n_1687),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1762),
.B(n_1675),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1769),
.Y(n_1834)
);

AND2x2_ASAP7_75t_SL g1835 ( 
.A(n_1768),
.B(n_1655),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1766),
.B(n_1672),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1751),
.B(n_1639),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1749),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1828),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1838),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1835),
.A2(n_1788),
.B1(n_1782),
.B2(n_1768),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_1836),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1805),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1833),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1805),
.B(n_1750),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1818),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1826),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1835),
.A2(n_1788),
.B1(n_1782),
.B2(n_1791),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1836),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1820),
.A2(n_1765),
.B(n_1799),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1838),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1821),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1814),
.B(n_1758),
.Y(n_1855)
);

OAI211xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1822),
.A2(n_1777),
.B(n_1801),
.C(n_1779),
.Y(n_1856)
);

OAI31xp33_ASAP7_75t_L g1857 ( 
.A1(n_1832),
.A2(n_1777),
.A3(n_1788),
.B(n_1643),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1822),
.A2(n_1801),
.B1(n_1788),
.B2(n_1779),
.C(n_1794),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1835),
.A2(n_1763),
.B1(n_1760),
.B2(n_1758),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1805),
.B(n_1810),
.Y(n_1861)
);

AOI21xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1832),
.A2(n_1657),
.B(n_1773),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1835),
.A2(n_1791),
.B1(n_1798),
.B2(n_1785),
.Y(n_1863)
);

OAI33xp33_ASAP7_75t_L g1864 ( 
.A1(n_1813),
.A2(n_1758),
.A3(n_1793),
.B1(n_1792),
.B2(n_1787),
.B3(n_1789),
.Y(n_1864)
);

NAND2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1811),
.B(n_1653),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1834),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1807),
.A2(n_1837),
.B1(n_1813),
.B2(n_1804),
.C(n_1814),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1834),
.Y(n_1868)
);

NAND2xp33_ASAP7_75t_R g1869 ( 
.A(n_1810),
.B(n_1796),
.Y(n_1869)
);

OAI31xp33_ASAP7_75t_L g1870 ( 
.A1(n_1807),
.A2(n_1659),
.A3(n_1644),
.B(n_1646),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1831),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1837),
.A2(n_1763),
.B1(n_1760),
.B2(n_1754),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1808),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1831),
.A2(n_1772),
.B1(n_1785),
.B2(n_1754),
.Y(n_1874)
);

OAI33xp33_ASAP7_75t_L g1875 ( 
.A1(n_1804),
.A2(n_1793),
.A3(n_1792),
.B1(n_1781),
.B2(n_1789),
.B3(n_1787),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1831),
.A2(n_1628),
.B1(n_1629),
.B2(n_1803),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_SL g1877 ( 
.A1(n_1824),
.A2(n_1776),
.B(n_1794),
.C(n_1781),
.Y(n_1877)
);

OAI33xp33_ASAP7_75t_L g1878 ( 
.A1(n_1823),
.A2(n_1795),
.A3(n_1802),
.B1(n_1797),
.B2(n_1770),
.B3(n_1775),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1820),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1811),
.A2(n_1791),
.B1(n_1798),
.B2(n_1785),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1816),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1817),
.B(n_1774),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1836),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1820),
.A2(n_1765),
.B(n_1799),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1816),
.Y(n_1885)
);

NOR2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1843),
.B(n_1824),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1881),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1847),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1853),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1843),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1881),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1867),
.B(n_1812),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1843),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1885),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1847),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1847),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1844),
.B(n_1806),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1857),
.B(n_1824),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1844),
.B(n_1806),
.Y(n_1900)
);

NOR2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1850),
.B(n_1883),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1873),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1851),
.A2(n_1820),
.B(n_1790),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1839),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1850),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1839),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1848),
.Y(n_1907)
);

OA21x2_ASAP7_75t_L g1908 ( 
.A1(n_1884),
.A2(n_1825),
.B(n_1827),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1874),
.B(n_1767),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1861),
.B(n_1806),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1854),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1854),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1859),
.A2(n_1791),
.B(n_1830),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1848),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1882),
.B(n_1827),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1868),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1868),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1840),
.Y(n_1919)
);

NOR3xp33_ASAP7_75t_L g1920 ( 
.A(n_1862),
.B(n_1741),
.C(n_1694),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1848),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1852),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1849),
.B(n_1829),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1848),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1866),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1863),
.A2(n_1798),
.B(n_1756),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1871),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1892),
.B(n_1862),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1892),
.B(n_1871),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1908),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1901),
.B(n_1861),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1899),
.B(n_1842),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1899),
.B(n_1842),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1901),
.B(n_1861),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1910),
.B(n_1927),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1894),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1910),
.B(n_1858),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1886),
.B(n_1861),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1894),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1887),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1886),
.B(n_1850),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1890),
.B(n_1883),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1911),
.B(n_1883),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1908),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1911),
.B(n_1846),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1927),
.B(n_1882),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1887),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1889),
.B(n_1858),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1908),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1919),
.B(n_1922),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1891),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1891),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1911),
.B(n_1846),
.Y(n_1953)
);

OR2x6_ASAP7_75t_L g1954 ( 
.A(n_1914),
.B(n_1759),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1889),
.B(n_1855),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1923),
.B(n_1872),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1923),
.B(n_1809),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1919),
.B(n_1809),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1893),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1893),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1913),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1926),
.B(n_1759),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1922),
.B(n_1809),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1894),
.B(n_1846),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1905),
.B(n_1846),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1925),
.B(n_1815),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1895),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1925),
.B(n_1815),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1905),
.B(n_1845),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1902),
.B(n_1815),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1905),
.B(n_1845),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1890),
.B(n_1879),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1895),
.Y(n_1973)
);

NOR3xp33_ASAP7_75t_L g1974 ( 
.A(n_1926),
.B(n_1877),
.C(n_1856),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1928),
.B(n_1902),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1974),
.B(n_1819),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1956),
.B(n_1860),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1935),
.B(n_1819),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1935),
.B(n_1904),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1936),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1940),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1931),
.B(n_1890),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1932),
.B(n_1864),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1954),
.A2(n_1841),
.B1(n_1880),
.B2(n_1909),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1950),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1940),
.Y(n_1986)
);

NAND2x1_ASAP7_75t_SL g1987 ( 
.A(n_1931),
.B(n_1909),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1947),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1947),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1934),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1936),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1951),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1929),
.B(n_1933),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1937),
.B(n_1819),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1951),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1952),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1952),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1957),
.B(n_1875),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1950),
.B(n_1904),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1939),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1946),
.B(n_1906),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1958),
.B(n_1920),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1963),
.B(n_1920),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1959),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1959),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1954),
.A2(n_1865),
.B1(n_1874),
.B2(n_1869),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1960),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1960),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1934),
.B(n_1898),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1938),
.B(n_1898),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1938),
.B(n_1898),
.Y(n_2011)
);

NOR2x1p5_ASAP7_75t_L g2012 ( 
.A(n_1975),
.B(n_1955),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1993),
.B(n_1979),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1982),
.B(n_1941),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1993),
.B(n_1939),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1981),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_L g2017 ( 
.A(n_1984),
.B(n_1961),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1980),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1982),
.B(n_1941),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1999),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1983),
.A2(n_1954),
.B1(n_1962),
.B2(n_1798),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1983),
.B(n_1948),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1980),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1985),
.B(n_1998),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1999),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1979),
.B(n_1946),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1998),
.A2(n_1954),
.B1(n_1962),
.B2(n_1965),
.Y(n_2028)
);

INVx1_ASAP7_75t_SL g2029 ( 
.A(n_1990),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1986),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1988),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1991),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1991),
.B(n_1961),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1989),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1992),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_2000),
.B(n_1978),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_2000),
.B(n_1967),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_2001),
.B(n_1967),
.Y(n_2039)
);

OA222x2_ASAP7_75t_L g2040 ( 
.A1(n_2015),
.A2(n_1954),
.B1(n_1962),
.B2(n_1987),
.C1(n_2003),
.C2(n_2002),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_SL g2041 ( 
.A1(n_2025),
.A2(n_2006),
.B(n_1976),
.Y(n_2041)
);

AOI222xp33_ASAP7_75t_L g2042 ( 
.A1(n_2017),
.A2(n_1977),
.B1(n_2010),
.B2(n_2011),
.C1(n_2007),
.C2(n_2005),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2033),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_2015),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2018),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2029),
.B(n_2010),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_2017),
.A2(n_1962),
.B(n_1995),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2021),
.A2(n_1962),
.B1(n_1994),
.B2(n_2011),
.Y(n_2048)
);

OAI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_2028),
.A2(n_2008),
.B1(n_2004),
.B2(n_1997),
.C(n_1996),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2018),
.Y(n_2050)
);

OAI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2022),
.A2(n_1870),
.B1(n_2001),
.B2(n_1876),
.C(n_1965),
.Y(n_2051)
);

AOI222xp33_ASAP7_75t_L g2052 ( 
.A1(n_2012),
.A2(n_1878),
.B1(n_1930),
.B2(n_1944),
.C1(n_1949),
.C2(n_1913),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2024),
.B(n_1970),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2024),
.B(n_1966),
.Y(n_2054)
);

INVxp67_ASAP7_75t_L g2055 ( 
.A(n_2013),
.Y(n_2055)
);

NAND4xp25_ASAP7_75t_SL g2056 ( 
.A(n_2014),
.B(n_1870),
.C(n_1943),
.D(n_1953),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_2013),
.B(n_1942),
.Y(n_2057)
);

O2A1O1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_2016),
.A2(n_1930),
.B(n_1944),
.C(n_1949),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2037),
.B(n_1968),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2014),
.B(n_1945),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2044),
.B(n_2020),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2055),
.B(n_2023),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2043),
.B(n_2023),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2045),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2046),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2060),
.B(n_2019),
.Y(n_2066)
);

NAND2x1p5_ASAP7_75t_L g2067 ( 
.A(n_2057),
.B(n_2034),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2042),
.B(n_2019),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2057),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_2041),
.B(n_2056),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2049),
.B(n_2037),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2050),
.B(n_2032),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_L g2073 ( 
.A(n_2047),
.B(n_2034),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2053),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2066),
.B(n_2032),
.Y(n_2075)
);

AOI221x1_ASAP7_75t_L g2076 ( 
.A1(n_2064),
.A2(n_2034),
.B1(n_2031),
.B2(n_2030),
.C(n_2035),
.Y(n_2076)
);

OR3x1_ASAP7_75t_L g2077 ( 
.A(n_2071),
.B(n_2026),
.C(n_2020),
.Y(n_2077)
);

OAI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2070),
.A2(n_2048),
.B(n_2051),
.Y(n_2078)
);

NAND4xp25_ASAP7_75t_L g2079 ( 
.A(n_2062),
.B(n_2059),
.C(n_2054),
.D(n_2052),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_SL g2080 ( 
.A(n_2067),
.B(n_2040),
.C(n_2059),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2068),
.B(n_2026),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_2073),
.A2(n_2036),
.B(n_2038),
.Y(n_2082)
);

NOR3xp33_ASAP7_75t_L g2083 ( 
.A(n_2065),
.B(n_2038),
.C(n_2027),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_L g2084 ( 
.A(n_2061),
.B(n_2027),
.C(n_2058),
.Y(n_2084)
);

OAI211xp5_ASAP7_75t_SL g2085 ( 
.A1(n_2069),
.A2(n_2039),
.B(n_1930),
.C(n_1949),
.Y(n_2085)
);

OAI222xp33_ASAP7_75t_L g2086 ( 
.A1(n_2067),
.A2(n_2039),
.B1(n_1944),
.B2(n_1972),
.C1(n_1942),
.C2(n_1971),
.Y(n_2086)
);

O2A1O1Ixp33_ASAP7_75t_SL g2087 ( 
.A1(n_2061),
.A2(n_1973),
.B(n_1917),
.C(n_1906),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_SL g2088 ( 
.A(n_2086),
.B(n_2063),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2080),
.A2(n_2072),
.B1(n_2074),
.B2(n_1942),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_R g2090 ( 
.A(n_2081),
.B(n_1969),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2075),
.B(n_1969),
.Y(n_2091)
);

OAI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_2079),
.A2(n_1942),
.B(n_1943),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_2083),
.B(n_1972),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2082),
.A2(n_1973),
.B(n_1972),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2090),
.B(n_2078),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2091),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2089),
.B(n_2084),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_2088),
.B(n_2085),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2092),
.B(n_2076),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2093),
.B(n_1945),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2094),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_L g2102 ( 
.A(n_2097),
.B(n_2077),
.Y(n_2102)
);

AOI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_2098),
.A2(n_2087),
.B(n_1972),
.C(n_1971),
.Y(n_2103)
);

OA22x2_ASAP7_75t_L g2104 ( 
.A1(n_2101),
.A2(n_1953),
.B1(n_1917),
.B2(n_1918),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2100),
.B(n_1913),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_2099),
.Y(n_2106)
);

AOI211x1_ASAP7_75t_SL g2107 ( 
.A1(n_2099),
.A2(n_1896),
.B(n_1897),
.C(n_1915),
.Y(n_2107)
);

NOR2x1_ASAP7_75t_L g2108 ( 
.A(n_2102),
.B(n_2095),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2106),
.B(n_2096),
.Y(n_2109)
);

NOR2x1_ASAP7_75t_L g2110 ( 
.A(n_2105),
.B(n_1913),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2108),
.B(n_2103),
.Y(n_2111)
);

OAI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_2111),
.A2(n_2109),
.B1(n_2110),
.B2(n_2107),
.C(n_2104),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_SL g2113 ( 
.A1(n_2112),
.A2(n_1912),
.B1(n_1918),
.B2(n_1916),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2112),
.A2(n_1916),
.B1(n_1912),
.B2(n_1896),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2113),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2114),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2115),
.A2(n_1916),
.B(n_1903),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_2116),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2118),
.A2(n_1897),
.B1(n_1896),
.B2(n_1915),
.Y(n_2119)
);

AOI221xp5_ASAP7_75t_L g2120 ( 
.A1(n_2119),
.A2(n_2117),
.B1(n_1897),
.B2(n_1896),
.C(n_1915),
.Y(n_2120)
);

AO21x2_ASAP7_75t_L g2121 ( 
.A1(n_2120),
.A2(n_1915),
.B(n_1897),
.Y(n_2121)
);

AOI22x1_ASAP7_75t_L g2122 ( 
.A1(n_2121),
.A2(n_1907),
.B1(n_1888),
.B2(n_1924),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_2122),
.A2(n_1900),
.B1(n_1924),
.B2(n_1921),
.Y(n_2123)
);

AOI211xp5_ASAP7_75t_L g2124 ( 
.A1(n_2123),
.A2(n_1853),
.B(n_1903),
.C(n_1888),
.Y(n_2124)
);


endmodule