module fake_jpeg_1693_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_63),
.B1(n_57),
.B2(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_48),
.B1(n_54),
.B2(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_75),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_54),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_66),
.B1(n_73),
.B2(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_46),
.B1(n_55),
.B2(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_46),
.B1(n_55),
.B2(n_53),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_91),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_62),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_1),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_44),
.B1(n_50),
.B2(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_50),
.B1(n_49),
.B2(n_3),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_2),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_98),
.B(n_104),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_96),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_92),
.B1(n_87),
.B2(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_5),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_1),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_21),
.B(n_36),
.C(n_35),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_22),
.B(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_17),
.C(n_34),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_26),
.C(n_25),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_122),
.B1(n_127),
.B2(n_6),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_123),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_37),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_6),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_24),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_94),
.B1(n_98),
.B2(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_109),
.B(n_23),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_122),
.B(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_109),
.B1(n_7),
.B2(n_8),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_9),
.C(n_10),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_123),
.C(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_117),
.C(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_121),
.B1(n_115),
.B2(n_13),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_144),
.A2(n_135),
.B1(n_130),
.B2(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_147),
.B1(n_142),
.B2(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_149),
.B1(n_133),
.B2(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_141),
.B1(n_121),
.B2(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_149),
.C(n_136),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_11),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_152),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_14),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_14),
.Y(n_156)
);


endmodule