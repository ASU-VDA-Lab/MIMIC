module real_jpeg_24065_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_63),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_37),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_46),
.B1(n_64),
.B2(n_65),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_69),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_81),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_9),
.A2(n_37),
.B1(n_40),
.B2(n_81),
.Y(n_132)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_37),
.B1(n_40),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_55),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_27),
.B1(n_37),
.B2(n_40),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_27),
.B1(n_64),
.B2(n_65),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_29),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_14),
.A2(n_42),
.B1(n_64),
.B2(n_65),
.Y(n_214)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_15),
.B(n_36),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_15),
.B(n_49),
.C(n_51),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_15),
.A2(n_37),
.B1(n_40),
.B2(n_111),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_106),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_111),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_15),
.B(n_64),
.C(n_76),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_15),
.A2(n_66),
.B(n_215),
.Y(n_245)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_16),
.Y(n_118)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_142),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_20),
.B(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_93),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_21),
.A2(n_22),
.B1(n_82),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_25),
.B(n_43),
.C(n_59),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_26),
.Y(n_95)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_30),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_30),
.A2(n_110),
.B(n_137),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_32),
.A2(n_37),
.B(n_110),
.C(n_112),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_33),
.B(n_34),
.C(n_40),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_35),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_35),
.B(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_37),
.B(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_41),
.Y(n_134)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_53),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_45),
.A2(n_47),
.B1(n_57),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_47),
.A2(n_53),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_49),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_49),
.B(n_224),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_54),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_104),
.B1(n_106),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_57),
.A2(n_105),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_72),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_60),
.B(n_72),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_113)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_65),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_65),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_68),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_70),
.B(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_66),
.A2(n_116),
.B1(n_118),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_66),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_66),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_73),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_73),
.A2(n_203),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_89),
.B1(n_90),
.B2(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_74),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_74),
.A2(n_90),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_78),
.A2(n_79),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_78),
.A2(n_153),
.B(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_78),
.B(n_111),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_82),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_92),
.Y(n_128)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_86),
.Y(n_230)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_90),
.B(n_154),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_93),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.C(n_107),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_94),
.B(n_102),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_111),
.CON(n_110),
.SN(n_110)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_107),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_111),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_114),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_118),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_139),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_172),
.B(n_263),
.C(n_268),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_166),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_156),
.C(n_159),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_145),
.A2(n_146),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_151),
.C(n_155),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_256),
.B(n_262),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_204),
.B(n_255),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_193),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_177),
.B(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.C(n_190),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B(n_184),
.Y(n_181)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_200),
.C(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_249),
.B(n_254),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_225),
.B(n_248),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_219),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_219),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_234),
.B(n_247),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_232),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_246),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);


endmodule