module fake_jpeg_5331_n_275 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_45),
.A2(n_48),
.B1(n_56),
.B2(n_33),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_36),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_21),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_1),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_34),
.B(n_36),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_2),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_24),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_23),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_71),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_73),
.Y(n_121)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_75),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_18),
.B1(n_34),
.B2(n_38),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_77),
.B1(n_102),
.B2(n_107),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_56),
.B1(n_48),
.B2(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_81),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_32),
.B(n_4),
.C(n_6),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_30),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_103),
.Y(n_126)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_16),
.Y(n_138)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_24),
.B1(n_33),
.B2(n_38),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_42),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_37),
.B(n_32),
.Y(n_124)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_33),
.B1(n_26),
.B2(n_30),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_108),
.A2(n_111),
.B1(n_3),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_41),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_115),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_41),
.B1(n_37),
.B2(n_29),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_114),
.A2(n_99),
.B1(n_73),
.B2(n_101),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_41),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_125),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_21),
.C(n_31),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_128),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_27),
.B1(n_37),
.B2(n_41),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_124),
.B1(n_141),
.B2(n_104),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_37),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_3),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_32),
.C(n_17),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_134),
.Y(n_169)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_67),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_3),
.C(n_6),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_32),
.B1(n_16),
.B2(n_15),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_145),
.Y(n_178)
);

NAND2x1_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_68),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_124),
.B(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_81),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_155),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_87),
.B1(n_88),
.B2(n_97),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_136),
.B1(n_127),
.B2(n_123),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_109),
.B(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_71),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_166),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_171),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_98),
.A3(n_101),
.B1(n_12),
.B2(n_13),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_130),
.B1(n_110),
.B2(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_179),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_166),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_129),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_186),
.B(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_119),
.C(n_118),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_143),
.C(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_198),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_163),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_202),
.B(n_211),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_144),
.B(n_167),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_192),
.B(n_183),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_157),
.C(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_142),
.C(n_160),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_120),
.B(n_9),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_156),
.C(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_198),
.C(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_7),
.B(n_10),
.C(n_11),
.D(n_13),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_15),
.C(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_147),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_190),
.B(n_177),
.Y(n_226)
);

AOI321xp33_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_201),
.A3(n_202),
.B1(n_190),
.B2(n_210),
.C(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_215),
.B1(n_204),
.B2(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_199),
.B1(n_213),
.B2(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_182),
.B1(n_212),
.B2(n_197),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_174),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_237),
.C(n_178),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_174),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_240),
.B(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_247),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_189),
.B1(n_182),
.B2(n_212),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_229),
.B(n_184),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_227),
.C(n_230),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_221),
.B(n_225),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_228),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_246),
.B1(n_245),
.B2(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_233),
.B1(n_225),
.B2(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_196),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_238),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_260),
.A2(n_223),
.B(n_147),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_256),
.A2(n_248),
.B1(n_239),
.B2(n_249),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_253),
.C(n_218),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_269),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_181),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_264),
.B(n_262),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_130),
.C(n_110),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_272),
.B(n_271),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_259),
.C(n_271),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_274),
.B(n_258),
.CI(n_273),
.CON(n_275),
.SN(n_275)
);


endmodule