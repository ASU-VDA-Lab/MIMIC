module fake_jpeg_14518_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_58),
.Y(n_183)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g207 ( 
.A(n_61),
.Y(n_207)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_66),
.B(n_72),
.Y(n_128)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_1),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_68),
.B(n_46),
.Y(n_191)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_70),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_19),
.B(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_80),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_87),
.Y(n_156)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_15),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_34),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_99),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_1),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_24),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_22),
.B1(n_46),
.B2(n_28),
.Y(n_141)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_35),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_107),
.B(n_108),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_35),
.B(n_45),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_118),
.Y(n_195)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_2),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_57),
.Y(n_120)
);

INVx5_ASAP7_75t_SL g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_20),
.Y(n_122)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_68),
.B(n_53),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_127),
.B(n_197),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_68),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_132),
.B(n_2),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_141),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_55),
.B1(n_23),
.B2(n_52),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_143),
.A2(n_157),
.B1(n_168),
.B2(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_72),
.B1(n_92),
.B2(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_145),
.A2(n_199),
.B1(n_191),
.B2(n_132),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_SL g147 ( 
.A(n_124),
.Y(n_147)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_74),
.A2(n_22),
.B1(n_46),
.B2(n_28),
.Y(n_157)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_61),
.Y(n_161)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_37),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_167),
.B(n_184),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_60),
.A2(n_55),
.B1(n_23),
.B2(n_52),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_81),
.B(n_43),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_43),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_187),
.B(n_192),
.Y(n_273)
);

NAND2x1_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_64),
.B(n_32),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_71),
.A2(n_30),
.B1(n_42),
.B2(n_37),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_75),
.B(n_42),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_97),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_77),
.A2(n_26),
.B1(n_53),
.B2(n_28),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_200),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_78),
.Y(n_203)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_86),
.B(n_79),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_210),
.B(n_214),
.Y(n_304)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_213),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_217),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_218),
.A2(n_264),
.B1(n_163),
.B2(n_189),
.Y(n_292)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_129),
.A2(n_179),
.B1(n_182),
.B2(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_221),
.A2(n_170),
.B1(n_158),
.B2(n_160),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_22),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_224),
.B(n_267),
.Y(n_299)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_225),
.Y(n_331)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_226),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_140),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_227),
.B(n_229),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_142),
.A2(n_198),
.B1(n_131),
.B2(n_169),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_230),
.A2(n_238),
.B1(n_266),
.B2(n_171),
.Y(n_302)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_129),
.A2(n_21),
.B(n_3),
.C(n_4),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_233),
.A2(n_207),
.B(n_151),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_152),
.A2(n_96),
.B1(n_93),
.B2(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_239),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_240),
.B(n_262),
.Y(n_324)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_242),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_243),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_207),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_127),
.B(n_3),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_249),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_156),
.B(n_13),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_250),
.C(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_4),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_4),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_253),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_254),
.A2(n_265),
.B1(n_272),
.B2(n_276),
.Y(n_315)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_149),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_195),
.B(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_139),
.B(n_6),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_149),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_157),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_183),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_271),
.Y(n_280)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_172),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_270),
.B(n_211),
.Y(n_329)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_166),
.A2(n_12),
.B1(n_190),
.B2(n_128),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_12),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_146),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_190),
.A2(n_12),
.B1(n_128),
.B2(n_186),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_204),
.B(n_154),
.C(n_137),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_133),
.C(n_170),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_189),
.B(n_174),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_230),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_260),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_281),
.B(n_284),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_291),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_286),
.B(n_326),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_292),
.A2(n_247),
.B1(n_250),
.B2(n_249),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g360 ( 
.A1(n_296),
.A2(n_213),
.B(n_263),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_220),
.B(n_133),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_300),
.B(n_312),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_308),
.B1(n_261),
.B2(n_243),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_244),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_313),
.C(n_322),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_307),
.A2(n_238),
.B1(n_256),
.B2(n_216),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_218),
.A2(n_151),
.B1(n_158),
.B2(n_160),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_244),
.A2(n_162),
.B(n_228),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_283),
.B(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_245),
.B(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_237),
.B(n_162),
.C(n_277),
.Y(n_313)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_237),
.B(n_246),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_269),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_234),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_328),
.A2(n_287),
.B(n_315),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_261),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_332),
.A2(n_337),
.B1(n_350),
.B2(n_355),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_336),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_233),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_257),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_338),
.B(n_344),
.Y(n_402)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_247),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_250),
.C(n_236),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_357),
.C(n_288),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_266),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_347),
.B(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_222),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_265),
.B1(n_271),
.B2(n_275),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_352),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_299),
.A2(n_215),
.B(n_263),
.Y(n_353)
);

HB1xp67_ASAP7_75t_SL g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_268),
.B1(n_259),
.B2(n_258),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_356),
.B(n_371),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_239),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_360),
.B1(n_367),
.B2(n_290),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_291),
.A2(n_262),
.B1(n_241),
.B2(n_223),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_359),
.A2(n_327),
.B1(n_280),
.B2(n_289),
.Y(n_377)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_311),
.Y(n_361)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_365),
.Y(n_394)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_315),
.A2(n_209),
.B1(n_248),
.B2(n_242),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_369),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_298),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_288),
.B(n_252),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_343),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_348),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_374),
.B(n_391),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_367),
.A2(n_304),
.B1(n_307),
.B2(n_321),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_377),
.A2(n_390),
.B1(n_395),
.B2(n_404),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_298),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_379),
.C(n_386),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_290),
.C(n_301),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_310),
.B(n_316),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_381),
.A2(n_310),
.B(n_318),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_290),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_338),
.B(n_282),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_332),
.A2(n_305),
.B1(n_255),
.B2(n_225),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_349),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_389),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_350),
.A2(n_219),
.B1(n_314),
.B2(n_231),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_317),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_397),
.A2(n_318),
.B(n_316),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_336),
.A2(n_282),
.B1(n_317),
.B2(n_325),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_383),
.A2(n_356),
.B1(n_337),
.B2(n_347),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_412),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_335),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_415),
.C(n_429),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_374),
.B(n_342),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_411),
.B(n_433),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_414),
.Y(n_447)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_383),
.A2(n_333),
.B1(n_359),
.B2(n_371),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_418),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_376),
.A2(n_342),
.B1(n_344),
.B2(n_366),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_426),
.Y(n_451)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_423),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_398),
.A2(n_340),
.B1(n_352),
.B2(n_370),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_430),
.B1(n_432),
.B2(n_400),
.Y(n_457)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_357),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

XOR2x1_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_346),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_428),
.B(n_379),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_353),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_368),
.B1(n_345),
.B2(n_363),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_431),
.A2(n_413),
.B(n_430),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_345),
.B1(n_365),
.B2(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_331),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_386),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_444),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_425),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_418),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_432),
.A2(n_384),
.B1(n_405),
.B2(n_393),
.Y(n_437)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_409),
.A2(n_382),
.B1(n_396),
.B2(n_402),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_456),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_415),
.C(n_407),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_435),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_428),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_449),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_396),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_452),
.A2(n_442),
.B(n_431),
.Y(n_476)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_453),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_382),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_458),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_409),
.A2(n_400),
.B1(n_393),
.B2(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_372),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_438),
.A2(n_408),
.B(n_412),
.Y(n_462)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_464),
.B(n_479),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_438),
.A2(n_451),
.B1(n_439),
.B2(n_424),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_456),
.B1(n_441),
.B2(n_443),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_427),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_478),
.Y(n_485)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_440),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_473),
.Y(n_493)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_459),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_385),
.Y(n_474)
);

AO221x1_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_394),
.B1(n_454),
.B2(n_447),
.C(n_426),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_476),
.A2(n_477),
.B1(n_463),
.B2(n_466),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_452),
.A2(n_408),
.B(n_433),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_480),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_372),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_377),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_405),
.B1(n_416),
.B2(n_421),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_404),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_468),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_466),
.A2(n_451),
.B1(n_434),
.B2(n_458),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_484),
.A2(n_475),
.B1(n_472),
.B2(n_462),
.Y(n_508)
);

BUFx24_ASAP7_75t_SL g486 ( 
.A(n_476),
.Y(n_486)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_446),
.C(n_448),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_492),
.C(n_497),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_444),
.C(n_455),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_467),
.A2(n_390),
.B1(n_443),
.B2(n_445),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_495),
.A2(n_465),
.B1(n_470),
.B2(n_460),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_420),
.C(n_414),
.Y(n_497)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_499),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_475),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_502),
.B(n_491),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_496),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_503),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_506),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_460),
.Y(n_506)
);

XNOR2x1_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_489),
.A2(n_423),
.B1(n_461),
.B2(n_381),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_510),
.A2(n_482),
.B1(n_487),
.B2(n_395),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_507),
.A2(n_483),
.B1(n_494),
.B2(n_495),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_512),
.A2(n_510),
.B1(n_507),
.B2(n_511),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_516),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_505),
.B(n_492),
.CI(n_484),
.CON(n_516),
.SN(n_516)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_517),
.A2(n_403),
.B1(n_397),
.B2(n_306),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_485),
.C(n_487),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_518),
.B(n_522),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_485),
.B(n_464),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_519),
.A2(n_508),
.B(n_509),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_461),
.C(n_401),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_524),
.A2(n_527),
.B(n_516),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_528),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_501),
.B(n_504),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_503),
.C(n_401),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_529),
.B(n_530),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_500),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_531),
.Y(n_532)
);

A2O1A1O1Ixp25_ASAP7_75t_L g533 ( 
.A1(n_523),
.A2(n_518),
.B(n_515),
.C(n_516),
.D(n_521),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_534),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_525),
.A2(n_515),
.B(n_513),
.Y(n_534)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_536),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_521),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_537),
.A2(n_529),
.B1(n_526),
.B2(n_403),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_540),
.A2(n_542),
.B(n_232),
.Y(n_545)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g541 ( 
.A1(n_535),
.A2(n_397),
.B(n_285),
.C(n_325),
.D(n_331),
.Y(n_541)
);

AOI321xp33_ASAP7_75t_SL g544 ( 
.A1(n_541),
.A2(n_295),
.A3(n_306),
.B1(n_285),
.B2(n_279),
.C(n_320),
.Y(n_544)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_538),
.C(n_532),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_543),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_545),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_540),
.C(n_279),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_547),
.B(n_295),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_226),
.B1(n_217),
.B2(n_235),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_235),
.Y(n_551)
);


endmodule