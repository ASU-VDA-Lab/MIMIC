module fake_aes_572_n_659 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_659);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_659;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_2), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_38), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_24), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_29), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_54), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_69), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_73), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_41), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_46), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_63), .Y(n_86) );
CKINVDCx14_ASAP7_75t_R g87 ( .A(n_47), .Y(n_87) );
INVx4_ASAP7_75t_R g88 ( .A(n_67), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_57), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_56), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_25), .Y(n_96) );
BUFx2_ASAP7_75t_L g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_32), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_72), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_27), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_51), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_30), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_17), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_22), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_61), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_31), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_5), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_18), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_62), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_43), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_103), .Y(n_122) );
INVx6_ASAP7_75t_L g123 ( .A(n_116), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_118), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_78), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_114), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_97), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g131 ( .A(n_77), .B(n_70), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_101), .B(n_0), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_87), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_102), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_84), .B(n_0), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_94), .B(n_66), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_114), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_76), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_79), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_76), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_104), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_112), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_113), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_105), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_80), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_106), .B(n_1), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_115), .B(n_2), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_108), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_80), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_109), .Y(n_159) );
INVxp67_ASAP7_75t_SL g160 ( .A(n_82), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_82), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_83), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_126), .B(n_127), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_126), .B(n_110), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_160), .B(n_121), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_127), .B(n_111), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_123), .Y(n_172) );
BUFx4f_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
BUFx12f_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_143), .B(n_120), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_122), .B(n_120), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_129), .B(n_119), .Y(n_178) );
INVx8_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
CKINVDCx8_ASAP7_75t_R g180 ( .A(n_135), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_123), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_135), .B(n_119), .Y(n_183) );
INVx6_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_146), .A2(n_117), .B1(n_100), .B2(n_99), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_162), .A2(n_92), .B1(n_100), .B2(n_99), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_139), .B(n_117), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_138), .B(n_98), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_98), .B1(n_96), .B2(n_95), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_134), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_140), .B(n_96), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_150), .B(n_95), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_150), .B(n_93), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_156), .B(n_93), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_123), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_152), .B(n_163), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_144), .A2(n_92), .B(n_91), .C(n_90), .Y(n_204) );
NAND3x1_ASAP7_75t_L g205 ( .A(n_154), .B(n_91), .C(n_90), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_156), .B(n_89), .C(n_86), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_163), .B(n_89), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_155), .B(n_86), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_162), .B(n_85), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_157), .B(n_137), .Y(n_213) );
OAI221xp5_ASAP7_75t_L g214 ( .A1(n_159), .A2(n_85), .B1(n_88), .B2(n_5), .C(n_6), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_159), .B(n_3), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_142), .B(n_3), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_203), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_168), .B(n_133), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_207), .Y(n_222) );
NOR2xp33_ASAP7_75t_R g223 ( .A(n_180), .B(n_124), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_212), .Y(n_224) );
NOR2xp33_ASAP7_75t_R g225 ( .A(n_180), .B(n_147), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_182), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_168), .B(n_153), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_168), .B(n_123), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_173), .A2(n_136), .B(n_125), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_177), .B(n_136), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_177), .B(n_125), .Y(n_233) );
NOR3xp33_ASAP7_75t_SL g234 ( .A(n_195), .B(n_4), .C(n_6), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_196), .B(n_163), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_190), .B(n_211), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_174), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_173), .A2(n_131), .B(n_163), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_173), .Y(n_241) );
OR2x2_ASAP7_75t_SL g242 ( .A(n_174), .B(n_4), .Y(n_242) );
NOR2x1p5_ASAP7_75t_L g243 ( .A(n_197), .B(n_7), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_190), .B(n_8), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_179), .Y(n_246) );
NAND3xp33_ASAP7_75t_SL g247 ( .A(n_194), .B(n_9), .C(n_10), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_165), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_211), .B(n_65), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_209), .B(n_9), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_166), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_214), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_197), .B(n_11), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_179), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_184), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_166), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_171), .B(n_12), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_181), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_181), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_197), .B(n_13), .Y(n_262) );
BUFx10_ASAP7_75t_L g263 ( .A(n_183), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_164), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_215), .B(n_13), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_181), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_179), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_184), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_215), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_205), .A2(n_26), .B(n_55), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_184), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_187), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_265), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_244), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_267), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_244), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_249), .A2(n_175), .B(n_193), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_267), .B(n_175), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_236), .B(n_178), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_227), .B(n_178), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_222), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_222), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_227), .B(n_198), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_255), .B(n_209), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_248), .B(n_200), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_237), .Y(n_296) );
BUFx8_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
CKINVDCx8_ASAP7_75t_R g298 ( .A(n_238), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_265), .A2(n_205), .B1(n_191), .B2(n_199), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_246), .B(n_206), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_278), .B(n_186), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_255), .B(n_176), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_277), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_224), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_250), .B(n_278), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
AND2x6_ASAP7_75t_L g309 ( .A(n_265), .B(n_185), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
NOR2x1_ASAP7_75t_SL g311 ( .A(n_256), .B(n_217), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_264), .B(n_167), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_249), .A2(n_208), .B(n_202), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_255), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_268), .B(n_169), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_240), .A2(n_208), .B(n_189), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_235), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_225), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_250), .B(n_213), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_277), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_260), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_223), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_257), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_262), .B(n_204), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_317), .B(n_262), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
OAI222xp33_ASAP7_75t_L g330 ( .A1(n_299), .A2(n_254), .B1(n_262), .B2(n_273), .C1(n_245), .C2(n_269), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_296), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_301), .A2(n_253), .B1(n_262), .B2(n_243), .Y(n_333) );
INVxp33_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
AOI21x1_ASAP7_75t_L g335 ( .A1(n_284), .A2(n_274), .B(n_229), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_309), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_286), .A2(n_254), .B1(n_247), .B2(n_230), .C(n_233), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_298), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
BUFx10_ASAP7_75t_L g343 ( .A(n_309), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_307), .B(n_253), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_318), .A2(n_274), .B(n_204), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_317), .B(n_269), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_310), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_326), .A2(n_253), .B1(n_243), .B2(n_252), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_315), .A2(n_253), .B1(n_259), .B2(n_256), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_293), .B(n_263), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_309), .A2(n_220), .B1(n_263), .B2(n_228), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_298), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_309), .B(n_263), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_309), .B(n_241), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_280), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_299), .B(n_234), .C(n_242), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_327), .B(n_307), .Y(n_359) );
AND2x6_ASAP7_75t_L g360 ( .A(n_336), .B(n_293), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_337), .A2(n_309), .B1(n_293), .B2(n_315), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_327), .A2(n_279), .B(n_289), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_337), .A2(n_287), .B1(n_292), .B2(n_316), .C(n_313), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_332), .A2(n_303), .B1(n_281), .B2(n_317), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_357), .A2(n_303), .B1(n_293), .B2(n_313), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g366 ( .A(n_333), .B(n_326), .C(n_321), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_357), .A2(n_326), .B1(n_317), .B2(n_289), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_326), .B1(n_302), .B2(n_263), .Y(n_369) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_290), .B(n_305), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_332), .B(n_281), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_356), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_329), .B(n_283), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_330), .A2(n_295), .B1(n_324), .B2(n_321), .C(n_288), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_300), .B(n_290), .C(n_306), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_335), .A2(n_318), .B(n_291), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_302), .B1(n_279), .B2(n_306), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_356), .Y(n_379) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_356), .B(n_283), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_328), .A2(n_302), .B1(n_282), .B2(n_288), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_344), .B(n_291), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_345), .B(n_297), .C(n_302), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_363), .B(n_338), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_365), .A2(n_352), .B(n_339), .C(n_353), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_375), .A2(n_328), .B1(n_351), .B2(n_352), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_384), .B(n_342), .Y(n_388) );
INVx5_ASAP7_75t_L g389 ( .A(n_360), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_382), .B(n_341), .Y(n_390) );
NAND2xp33_ASAP7_75t_SL g391 ( .A(n_381), .B(n_342), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_361), .A2(n_341), .B(n_347), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_373), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_361), .A2(n_328), .B1(n_342), .B2(n_336), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_380), .B(n_345), .C(n_350), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_366), .A2(n_330), .B1(n_347), .B2(n_349), .C(n_305), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_369), .A2(n_349), .B1(n_350), .B2(n_319), .C(n_351), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_358), .Y(n_398) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_371), .A2(n_202), .B(n_354), .C(n_340), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_367), .A2(n_351), .B1(n_328), .B2(n_342), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_383), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_383), .A2(n_319), .B1(n_282), .B2(n_213), .C(n_314), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_382), .B(n_282), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_359), .A2(n_354), .B1(n_346), .B2(n_285), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_345), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_364), .A2(n_285), .B1(n_346), .B2(n_241), .C(n_340), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_372), .B(n_345), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_340), .B1(n_355), .B2(n_270), .C(n_285), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_379), .B(n_340), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_360), .A2(n_297), .B1(n_355), .B2(n_331), .Y(n_412) );
AOI33xp33_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_188), .A3(n_216), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_346), .B1(n_355), .B2(n_322), .Y(n_414) );
NAND2xp33_ASAP7_75t_R g415 ( .A(n_374), .B(n_345), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_379), .A2(n_380), .B1(n_368), .B2(n_346), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_368), .Y(n_417) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_403), .B(n_343), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_406), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_406), .B(n_370), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_408), .B(n_370), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_393), .B(n_401), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_408), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_401), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_370), .Y(n_425) );
OAI21xp33_ASAP7_75t_SL g426 ( .A1(n_413), .A2(n_362), .B(n_346), .Y(n_426) );
INVxp33_ASAP7_75t_L g427 ( .A(n_403), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_392), .B(n_377), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_391), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_385), .B(n_377), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_387), .A2(n_346), .B1(n_304), .B2(n_322), .C(n_377), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_411), .B(n_377), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_394), .A2(n_360), .B1(n_355), .B2(n_343), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_411), .B(n_360), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
AND4x1_ASAP7_75t_SL g441 ( .A(n_387), .B(n_331), .C(n_343), .D(n_297), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_395), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_386), .B(n_331), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_396), .B(n_188), .C(n_216), .D(n_19), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_415), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_390), .B(n_360), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_360), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_399), .B(n_297), .C(n_304), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_394), .B(n_360), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_405), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_322), .B(n_325), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_395), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_404), .A2(n_323), .B(n_325), .Y(n_455) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_407), .B(n_172), .C(n_201), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_388), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_389), .B(n_14), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_389), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_389), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_389), .B(n_15), .Y(n_464) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_444), .B(n_414), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_426), .A2(n_409), .B(n_400), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_19), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_451), .B(n_397), .Y(n_468) );
NAND4xp75_ASAP7_75t_L g469 ( .A(n_443), .B(n_402), .C(n_343), .D(n_22), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_427), .B(n_20), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
OR2x4_ASAP7_75t_L g473 ( .A(n_462), .B(n_20), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_430), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_459), .B(n_21), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_459), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_430), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_420), .B(n_21), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_419), .B(n_423), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_420), .B(n_23), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
NOR4xp25_ASAP7_75t_SL g485 ( .A(n_432), .B(n_311), .C(n_33), .D(n_34), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_420), .B(n_28), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_419), .B(n_311), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_429), .B(n_323), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_461), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_423), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_421), .B(n_325), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_421), .B(n_325), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_421), .B(n_294), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_444), .B(n_426), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_461), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_450), .B(n_44), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_448), .B(n_312), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_450), .B(n_45), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_450), .B(n_49), .Y(n_500) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_449), .B(n_312), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_461), .B(n_50), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_425), .B(n_52), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_430), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_447), .B(n_312), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_441), .B(n_172), .C(n_201), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_464), .A2(n_312), .B1(n_294), .B2(n_226), .Y(n_507) );
BUFx12f_ASAP7_75t_L g508 ( .A(n_464), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_445), .A2(n_270), .B1(n_201), .B2(n_294), .C(n_226), .Y(n_509) );
NAND2xp33_ASAP7_75t_R g510 ( .A(n_458), .B(n_64), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_463), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_431), .B(n_226), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_435), .Y(n_513) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_457), .B(n_294), .C(n_323), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_448), .B(n_447), .Y(n_515) );
INVx3_ASAP7_75t_SL g516 ( .A(n_418), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_425), .B(n_226), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_435), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_425), .B(n_231), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_470), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_480), .B(n_448), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_477), .B(n_431), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
NAND5xp2_ASAP7_75t_L g525 ( .A(n_495), .B(n_432), .C(n_437), .D(n_464), .E(n_446), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g526 ( .A1(n_495), .A2(n_446), .B(n_457), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_465), .B(n_454), .C(n_453), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_510), .A2(n_429), .B1(n_462), .B2(n_449), .Y(n_529) );
INVxp33_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_483), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_481), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_510), .A2(n_445), .B1(n_438), .B2(n_418), .Y(n_535) );
OAI22xp33_ASAP7_75t_SL g536 ( .A1(n_467), .A2(n_463), .B1(n_454), .B2(n_458), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_468), .B(n_436), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_484), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_489), .A2(n_463), .B(n_460), .C(n_458), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_466), .A2(n_452), .B1(n_442), .B2(n_453), .C(n_460), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_471), .A2(n_433), .B1(n_434), .B2(n_438), .C1(n_442), .C2(n_453), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_501), .A2(n_455), .B(n_460), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g544 ( .A1(n_502), .A2(n_418), .A3(n_452), .B(n_458), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_516), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_485), .A2(n_455), .B(n_435), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_469), .A2(n_456), .B(n_442), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_479), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_516), .Y(n_550) );
XNOR2x1_ASAP7_75t_L g551 ( .A(n_482), .B(n_438), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_491), .B(n_515), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_504), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_513), .Y(n_554) );
OAI21xp5_ASAP7_75t_SL g555 ( .A1(n_502), .A2(n_441), .B(n_456), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_479), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_475), .A2(n_433), .B1(n_434), .B2(n_436), .C(n_428), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_508), .A2(n_436), .B1(n_428), .B2(n_440), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_517), .B(n_440), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_482), .A2(n_440), .B(n_231), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_518), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_514), .A2(n_231), .B(n_277), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_486), .A2(n_231), .B(n_275), .C(n_232), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_486), .A2(n_277), .B(n_232), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_494), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_517), .B(n_232), .Y(n_568) );
AO22x1_ASAP7_75t_L g569 ( .A1(n_511), .A2(n_277), .B1(n_232), .B2(n_275), .Y(n_569) );
XNOR2x2_ASAP7_75t_SL g570 ( .A(n_529), .B(n_473), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_524), .Y(n_571) );
INVx4_ASAP7_75t_L g572 ( .A(n_569), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_536), .B(n_511), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_545), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g575 ( .A(n_550), .B(n_500), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_552), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_528), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_520), .B(n_496), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_538), .B(n_519), .Y(n_579) );
AO22x2_ASAP7_75t_L g580 ( .A1(n_521), .A2(n_490), .B1(n_518), .B2(n_500), .Y(n_580) );
NOR4xp25_ASAP7_75t_SL g581 ( .A(n_526), .B(n_473), .C(n_508), .D(n_509), .Y(n_581) );
NOR4xp25_ASAP7_75t_SL g582 ( .A(n_555), .B(n_497), .C(n_499), .D(n_503), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_557), .B(n_519), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_551), .A2(n_497), .B1(n_499), .B2(n_503), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_534), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_520), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_540), .A2(n_487), .B(n_498), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_542), .B(n_512), .Y(n_588) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_558), .B(n_512), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_559), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_525), .B(n_505), .Y(n_591) );
XOR2xp5_ASAP7_75t_L g592 ( .A(n_551), .B(n_507), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_565), .B(n_567), .Y(n_593) );
NAND2xp33_ASAP7_75t_R g594 ( .A(n_564), .B(n_506), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_530), .B(n_260), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_531), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_527), .B(n_257), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_522), .B(n_221), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_523), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_544), .A2(n_275), .B(n_239), .Y(n_603) );
INVxp33_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_558), .B(n_221), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_586), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_585), .Y(n_608) );
AO22x2_ASAP7_75t_L g609 ( .A1(n_573), .A2(n_566), .B1(n_548), .B2(n_553), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_591), .A2(n_535), .B1(n_547), .B2(n_560), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_573), .A2(n_603), .B(n_591), .C(n_588), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_600), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g613 ( .A1(n_580), .A2(n_540), .A3(n_541), .B(n_563), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g614 ( .A1(n_584), .A2(n_543), .B1(n_568), .B2(n_554), .C1(n_546), .C2(n_556), .Y(n_614) );
AO22x2_ASAP7_75t_L g615 ( .A1(n_576), .A2(n_561), .B1(n_556), .B2(n_549), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_594), .A2(n_561), .B1(n_549), .B2(n_537), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_571), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_589), .A2(n_562), .B(n_537), .C(n_532), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_572), .A2(n_277), .B(n_239), .Y(n_619) );
BUFx8_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_577), .Y(n_621) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_582), .A2(n_275), .B(n_239), .C(n_251), .Y(n_622) );
OR3x1_ASAP7_75t_L g623 ( .A(n_570), .B(n_260), .C(n_251), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_572), .B(n_221), .C(n_251), .Y(n_624) );
AOI32xp33_ASAP7_75t_L g625 ( .A1(n_572), .A2(n_258), .A3(n_261), .B1(n_266), .B2(n_271), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_601), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_601), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_609), .B(n_580), .Y(n_628) );
OAI322xp33_ASAP7_75t_L g629 ( .A1(n_610), .A2(n_583), .A3(n_602), .B1(n_592), .B2(n_593), .C1(n_590), .C2(n_575), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_627), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_609), .A2(n_581), .B(n_580), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_623), .A2(n_604), .B1(n_579), .B2(n_578), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_611), .A2(n_604), .B1(n_597), .B2(n_596), .C(n_587), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_606), .B(n_598), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_613), .A2(n_594), .B1(n_595), .B2(n_605), .C(n_266), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_608), .B(n_595), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_614), .A2(n_258), .B(n_261), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_607), .B(n_258), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_617), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_610), .A2(n_261), .B1(n_266), .B2(n_271), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_622), .B(n_271), .C(n_272), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_618), .A2(n_272), .B(n_276), .C(n_260), .Y(n_643) );
NOR3xp33_ASAP7_75t_SL g644 ( .A(n_619), .B(n_260), .C(n_276), .Y(n_644) );
AOI211x1_ASAP7_75t_L g645 ( .A1(n_621), .A2(n_260), .B(n_272), .C(n_276), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_624), .A2(n_620), .B1(n_626), .B2(n_615), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_615), .A2(n_625), .B(n_616), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_628), .A2(n_646), .B1(n_636), .B2(n_631), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_635), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_620), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_630), .Y(n_651) );
NOR4xp25_ASAP7_75t_L g652 ( .A(n_648), .B(n_629), .C(n_634), .D(n_638), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_651), .B(n_647), .C(n_632), .Y(n_653) );
OR3x1_ASAP7_75t_L g654 ( .A(n_649), .B(n_633), .C(n_640), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_653), .A2(n_649), .B1(n_650), .B2(n_637), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_652), .A2(n_643), .B(n_641), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_655), .A2(n_654), .B1(n_616), .B2(n_639), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_656), .B1(n_642), .B2(n_639), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_645), .B(n_644), .Y(n_659) );
endmodule