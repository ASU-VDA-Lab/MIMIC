module real_aes_8309_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_1), .A2(n_164), .B(n_167), .C(n_247), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_2), .A2(n_193), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g494 ( .A(n_3), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_4), .B(n_223), .Y(n_222) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_5), .A2(n_193), .B(n_478), .Y(n_477) );
AND2x6_ASAP7_75t_L g164 ( .A(n_6), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g260 ( .A(n_7), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_8), .B(n_41), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_8), .B(n_41), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_9), .A2(n_192), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_10), .B(n_176), .Y(n_249) );
INVx1_ASAP7_75t_L g482 ( .A(n_11), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_12), .B(n_217), .Y(n_517) );
INVx1_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
INVx1_ASAP7_75t_L g529 ( .A(n_14), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_15), .A2(n_78), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_15), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_16), .A2(n_201), .B(n_282), .C(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_17), .B(n_223), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_18), .B(n_460), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_19), .B(n_193), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_20), .B(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_21), .A2(n_217), .B(n_268), .C(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_22), .B(n_223), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_23), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_24), .A2(n_203), .B(n_284), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_25), .B(n_176), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g158 ( .A(n_26), .Y(n_158) );
INVx1_ASAP7_75t_L g230 ( .A(n_27), .Y(n_230) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_28), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_29), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_30), .B(n_176), .Y(n_495) );
INVx1_ASAP7_75t_L g199 ( .A(n_31), .Y(n_199) );
INVx1_ASAP7_75t_L g472 ( .A(n_32), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_33), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_33), .Y(n_134) );
INVx2_ASAP7_75t_L g162 ( .A(n_34), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_35), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_36), .A2(n_217), .B(n_218), .C(n_220), .Y(n_216) );
INVxp67_ASAP7_75t_L g202 ( .A(n_37), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g215 ( .A(n_38), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_39), .A2(n_167), .B(n_229), .C(n_233), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_40), .A2(n_164), .B(n_167), .C(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g471 ( .A(n_42), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_43), .A2(n_178), .B(n_258), .C(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_44), .B(n_176), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_45), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_46), .Y(n_195) );
INVx1_ASAP7_75t_L g266 ( .A(n_47), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_48), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_49), .A2(n_58), .B1(n_742), .B2(n_743), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_49), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_50), .B(n_193), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_51), .A2(n_167), .B1(n_270), .B2(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_52), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_53), .Y(n_491) );
CKINVDCx14_ASAP7_75t_R g256 ( .A(n_54), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_55), .A2(n_220), .B(n_258), .C(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_56), .Y(n_541) );
INVx1_ASAP7_75t_L g479 ( .A(n_57), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_58), .Y(n_743) );
INVx1_ASAP7_75t_L g165 ( .A(n_59), .Y(n_165) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
INVx1_ASAP7_75t_SL g219 ( .A(n_61), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_62), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_63), .A2(n_741), .B1(n_744), .B2(n_745), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_63), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_64), .B(n_223), .Y(n_272) );
INVx1_ASAP7_75t_L g171 ( .A(n_65), .Y(n_171) );
AOI222xp33_ASAP7_75t_SL g131 ( .A1(n_66), .A2(n_132), .B1(n_133), .B2(n_139), .C1(n_732), .C2(n_734), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_SL g459 ( .A1(n_67), .A2(n_220), .B(n_460), .C(n_461), .Y(n_459) );
INVxp67_ASAP7_75t_L g462 ( .A(n_68), .Y(n_462) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_70), .A2(n_193), .B(n_255), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_71), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_72), .A2(n_193), .B(n_279), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_73), .Y(n_475) );
INVx1_ASAP7_75t_L g535 ( .A(n_74), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_75), .A2(n_192), .B(n_194), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_76), .Y(n_227) );
INVx1_ASAP7_75t_L g280 ( .A(n_77), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_78), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_79), .A2(n_164), .B(n_167), .C(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_80), .A2(n_193), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g283 ( .A(n_81), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_82), .B(n_200), .Y(n_506) );
INVx2_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx1_ASAP7_75t_L g248 ( .A(n_84), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_85), .B(n_460), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_86), .A2(n_164), .B(n_167), .C(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g126 ( .A(n_87), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g446 ( .A(n_87), .B(n_128), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_88), .A2(n_167), .B(n_170), .C(n_180), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_89), .B(n_185), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_90), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_91), .A2(n_164), .B(n_167), .C(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_92), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_93), .A2(n_104), .B1(n_117), .B2(n_747), .Y(n_103) );
INVx1_ASAP7_75t_L g458 ( .A(n_94), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_95), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_96), .B(n_200), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_98), .B(n_151), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_99), .B(n_151), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g269 ( .A(n_101), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_102), .A2(n_193), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g748 ( .A(n_107), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g128 ( .A(n_112), .B(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g731 ( .A(n_113), .B(n_128), .Y(n_731) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_113), .B(n_127), .Y(n_736) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_131), .B1(n_737), .B2(n_738), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g737 ( .A(n_122), .Y(n_737) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_124), .A2(n_739), .B(n_746), .Y(n_738) );
NOR2xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_130), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_126), .Y(n_746) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_446), .B1(n_447), .B2(n_729), .Y(n_139) );
INVx2_ASAP7_75t_L g733 ( .A(n_140), .Y(n_733) );
XOR2xp5_ASAP7_75t_L g739 ( .A(n_140), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_380), .Y(n_140) );
NAND5xp2_ASAP7_75t_L g141 ( .A(n_142), .B(n_309), .C(n_339), .D(n_360), .E(n_366), .Y(n_141) );
AOI221xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_239), .B1(n_273), .B2(n_275), .C(n_286), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_236), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_208), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_SL g360 ( .A1(n_147), .A2(n_224), .B(n_361), .C(n_364), .Y(n_360) );
AND2x2_ASAP7_75t_L g430 ( .A(n_147), .B(n_225), .Y(n_430) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_186), .Y(n_147) );
AND2x2_ASAP7_75t_L g288 ( .A(n_148), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g292 ( .A(n_148), .B(n_289), .Y(n_292) );
OR2x2_ASAP7_75t_L g318 ( .A(n_148), .B(n_225), .Y(n_318) );
AND2x2_ASAP7_75t_L g320 ( .A(n_148), .B(n_211), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_148), .B(n_210), .Y(n_338) );
INVx1_ASAP7_75t_L g371 ( .A(n_148), .Y(n_371) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
BUFx2_ASAP7_75t_L g238 ( .A(n_149), .Y(n_238) );
AND2x2_ASAP7_75t_L g274 ( .A(n_149), .B(n_211), .Y(n_274) );
AND2x2_ASAP7_75t_L g427 ( .A(n_149), .B(n_225), .Y(n_427) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_157), .B(n_182), .Y(n_149) );
INVx3_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_150), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_150), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g508 ( .A(n_150), .B(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_151), .A2(n_456), .B(n_463), .Y(n_455) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_153), .B(n_154), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_166), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_159), .A2(n_185), .B(n_227), .C(n_228), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_159), .A2(n_245), .B(n_246), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_159), .A2(n_181), .B1(n_469), .B2(n_473), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_159), .A2(n_491), .B(n_492), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_159), .A2(n_535), .B(n_536), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AND2x4_ASAP7_75t_L g193 ( .A(n_160), .B(n_164), .Y(n_193) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
INVx1_ASAP7_75t_L g271 ( .A(n_162), .Y(n_271) );
INVx1_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
INVx3_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
INVx1_ASAP7_75t_L g460 ( .A(n_163), .Y(n_460) );
INVx4_ASAP7_75t_SL g181 ( .A(n_164), .Y(n_181) );
BUFx3_ASAP7_75t_L g233 ( .A(n_164), .Y(n_233) );
INVx5_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
AND2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
BUFx3_ASAP7_75t_L g179 ( .A(n_168), .Y(n_179) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_175), .C(n_177), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_172), .A2(n_177), .B(n_248), .C(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_173), .A2(n_174), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g203 ( .A(n_174), .Y(n_203) );
INVx4_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
INVx2_ASAP7_75t_L g258 ( .A(n_176), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_177), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_177), .A2(n_538), .B(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g284 ( .A(n_179), .Y(n_284) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_181), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_196), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_181), .A2(n_196), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_181), .A2(n_196), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_181), .A2(n_196), .B(n_280), .C(n_281), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_181), .A2(n_196), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_181), .A2(n_196), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_181), .A2(n_196), .B(n_526), .C(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_184), .A2(n_513), .B(n_520), .Y(n_512) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_254), .B(n_261), .Y(n_253) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_185), .A2(n_524), .B(n_530), .Y(n_523) );
AND2x2_ASAP7_75t_L g308 ( .A(n_186), .B(n_209), .Y(n_308) );
OR2x2_ASAP7_75t_L g312 ( .A(n_186), .B(n_225), .Y(n_312) );
AND2x2_ASAP7_75t_L g337 ( .A(n_186), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g384 ( .A(n_186), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_186), .B(n_346), .Y(n_432) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B(n_205), .Y(n_186) );
INVx1_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_187), .A2(n_534), .B(n_540), .Y(n_533) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_SL g502 ( .A1(n_188), .A2(n_503), .B(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_189), .A2(n_468), .B(n_474), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_189), .B(n_475), .Y(n_474) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_189), .A2(n_490), .B(n_497), .Y(n_489) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_191), .A2(n_206), .B(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_198), .B(n_204), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B1(n_202), .B2(n_203), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_200), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_200), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_201), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_201), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_201), .B(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_203), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_203), .B(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_203), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g232 ( .A(n_204), .Y(n_232) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OAI322xp33_ASAP7_75t_L g433 ( .A1(n_208), .A2(n_369), .A3(n_392), .B1(n_413), .B2(n_434), .C1(n_436), .C2(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_209), .B(n_289), .Y(n_436) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_224), .Y(n_209) );
AND2x2_ASAP7_75t_L g237 ( .A(n_210), .B(n_238), .Y(n_237) );
AND2x4_ASAP7_75t_L g305 ( .A(n_210), .B(n_225), .Y(n_305) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g346 ( .A(n_211), .B(n_225), .Y(n_346) );
AND2x2_ASAP7_75t_L g390 ( .A(n_211), .B(n_224), .Y(n_390) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_222), .Y(n_211) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_212), .A2(n_264), .B(n_272), .Y(n_263) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_212), .A2(n_278), .B(n_285), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_217), .B(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_221), .Y(n_518) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_223), .A2(n_477), .B(n_483), .Y(n_476) );
AND2x2_ASAP7_75t_L g273 ( .A(n_224), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g291 ( .A(n_224), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_224), .B(n_320), .Y(n_444) );
INVx3_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g236 ( .A(n_225), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_225), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g358 ( .A(n_225), .B(n_289), .Y(n_358) );
AND2x2_ASAP7_75t_L g385 ( .A(n_225), .B(n_320), .Y(n_385) );
OR2x2_ASAP7_75t_L g441 ( .A(n_225), .B(n_292), .Y(n_441) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_234), .Y(n_225) );
INVx1_ASAP7_75t_SL g327 ( .A(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_237), .B(n_358), .Y(n_359) );
AND2x2_ASAP7_75t_L g393 ( .A(n_237), .B(n_383), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_237), .B(n_316), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_237), .B(n_438), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_239), .A2(n_273), .A3(n_412), .B(n_414), .Y(n_411) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_252), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_240), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g394 ( .A(n_240), .B(n_329), .Y(n_394) );
OR2x2_ASAP7_75t_L g401 ( .A(n_240), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g413 ( .A(n_240), .B(n_302), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g347 ( .A(n_241), .B(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g275 ( .A(n_242), .B(n_276), .Y(n_275) );
INVx4_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
AND2x2_ASAP7_75t_L g333 ( .A(n_242), .B(n_277), .Y(n_333) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_250), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_243), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_243), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_243), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g332 ( .A(n_252), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g402 ( .A(n_252), .Y(n_402) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_262), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_253), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_263), .Y(n_302) );
INVx2_ASAP7_75t_L g322 ( .A(n_253), .Y(n_322) );
AND2x2_ASAP7_75t_L g336 ( .A(n_253), .B(n_263), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_299), .Y(n_343) );
BUFx3_ASAP7_75t_L g353 ( .A(n_253), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_253), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_296), .Y(n_306) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_263), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_263), .Y(n_330) );
INVx2_ASAP7_75t_L g496 ( .A(n_270), .Y(n_496) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_SL g313 ( .A(n_274), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_274), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_274), .B(n_383), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_275), .B(n_353), .Y(n_406) );
INVx1_ASAP7_75t_SL g440 ( .A(n_275), .Y(n_440) );
INVx1_ASAP7_75t_SL g348 ( .A(n_276), .Y(n_348) );
INVx1_ASAP7_75t_SL g299 ( .A(n_277), .Y(n_299) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
OR2x2_ASAP7_75t_L g321 ( .A(n_277), .B(n_296), .Y(n_321) );
AND2x2_ASAP7_75t_L g335 ( .A(n_277), .B(n_296), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_277), .B(n_325), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B(n_293), .C(n_304), .Y(n_286) );
AOI31xp33_ASAP7_75t_L g403 ( .A1(n_287), .A2(n_404), .A3(n_405), .B(n_406), .Y(n_403) );
AND2x2_ASAP7_75t_L g376 ( .A(n_288), .B(n_305), .Y(n_376) );
BUFx3_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_289), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g352 ( .A(n_289), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_289), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g307 ( .A(n_292), .Y(n_307) );
OAI222xp33_ASAP7_75t_L g416 ( .A1(n_292), .A2(n_417), .B1(n_420), .B2(n_421), .C1(n_422), .C2(n_423), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_300), .Y(n_293) );
INVx1_ASAP7_75t_L g422 ( .A(n_294), .Y(n_422) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_296), .B(n_299), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_296), .B(n_322), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_296), .B(n_297), .Y(n_392) );
INVx1_ASAP7_75t_L g443 ( .A(n_296), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_297), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g445 ( .A(n_297), .Y(n_445) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g325 ( .A(n_298), .Y(n_325) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
AOI32xp33_ASAP7_75t_L g304 ( .A1(n_300), .A2(n_305), .A3(n_306), .B1(n_307), .B2(n_308), .Y(n_304) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_302), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g379 ( .A(n_302), .Y(n_379) );
OR2x2_ASAP7_75t_L g420 ( .A(n_302), .B(n_321), .Y(n_420) );
INVx1_ASAP7_75t_L g356 ( .A(n_303), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_305), .B(n_316), .Y(n_341) );
INVx3_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
AOI322xp5_ASAP7_75t_L g366 ( .A1(n_305), .A2(n_350), .A3(n_367), .B1(n_369), .B2(n_372), .C1(n_376), .C2(n_377), .Y(n_366) );
AND2x2_ASAP7_75t_L g342 ( .A(n_306), .B(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g419 ( .A(n_306), .Y(n_419) );
A2O1A1O1Ixp25_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_314), .C(n_322), .D(n_323), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_310), .B(n_353), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_312), .A2(n_324), .B1(n_327), .B2(n_328), .C(n_331), .Y(n_323) );
INVx1_ASAP7_75t_SL g438 ( .A(n_312), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_319), .B(n_321), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_316), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_318), .A2(n_402), .B1(n_409), .B2(n_410), .C(n_411), .Y(n_408) );
OAI222xp33_ASAP7_75t_L g439 ( .A1(n_319), .A2(n_440), .B1(n_441), .B2(n_442), .C1(n_444), .C2(n_445), .Y(n_439) );
AND2x2_ASAP7_75t_L g397 ( .A(n_320), .B(n_383), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_320), .A2(n_335), .B(n_382), .Y(n_409) );
INVx1_ASAP7_75t_L g423 ( .A(n_320), .Y(n_423) );
INVx2_ASAP7_75t_SL g326 ( .A(n_321), .Y(n_326) );
AND2x2_ASAP7_75t_L g329 ( .A(n_322), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_SL g363 ( .A(n_325), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_325), .B(n_335), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_326), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_326), .B(n_336), .Y(n_365) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_337), .Y(n_331) );
INVx1_ASAP7_75t_SL g349 ( .A(n_333), .Y(n_349) );
AND2x2_ASAP7_75t_L g396 ( .A(n_333), .B(n_379), .Y(n_396) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x2_ASAP7_75t_L g435 ( .A(n_335), .B(n_353), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_336), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g421 ( .A(n_337), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_344), .B2(n_351), .C(n_354), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_349), .B2(n_350), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_348), .A2(n_355), .B1(n_357), .B2(n_359), .Y(n_354) );
OR2x2_ASAP7_75t_L g425 ( .A(n_349), .B(n_353), .Y(n_425) );
OR2x2_ASAP7_75t_L g428 ( .A(n_349), .B(n_363), .Y(n_428) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_425), .B1(n_426), .B2(n_428), .C(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_395), .C(n_407), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_386), .B1(n_388), .B2(n_391), .C1(n_393), .C2(n_394), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_383), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g410 ( .A(n_396), .Y(n_410) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_400), .A2(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NOR5xp2_ASAP7_75t_L g407 ( .A(n_408), .B(n_416), .C(n_424), .D(n_433), .E(n_439), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_446), .A2(n_448), .B1(n_729), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_449), .B(n_666), .Y(n_448) );
NOR4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_596), .C(n_627), .D(n_646), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_554), .C(n_569), .D(n_587), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_499), .B1(n_531), .B2(n_542), .C1(n_547), .C2(n_549), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_484), .Y(n_452) );
INVx1_ASAP7_75t_L g610 ( .A(n_453), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_464), .Y(n_453) );
AND2x2_ASAP7_75t_L g485 ( .A(n_454), .B(n_476), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_454), .B(n_488), .Y(n_639) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g546 ( .A(n_455), .B(n_466), .Y(n_546) );
AND2x2_ASAP7_75t_L g555 ( .A(n_455), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g581 ( .A(n_455), .Y(n_581) );
AND2x2_ASAP7_75t_L g602 ( .A(n_455), .B(n_466), .Y(n_602) );
BUFx2_ASAP7_75t_L g625 ( .A(n_455), .Y(n_625) );
AND2x2_ASAP7_75t_L g649 ( .A(n_455), .B(n_467), .Y(n_649) );
AND2x2_ASAP7_75t_L g713 ( .A(n_455), .B(n_476), .Y(n_713) );
AND2x2_ASAP7_75t_L g614 ( .A(n_464), .B(n_545), .Y(n_614) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_465), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
OR2x2_ASAP7_75t_L g574 ( .A(n_466), .B(n_489), .Y(n_574) );
AND2x2_ASAP7_75t_L g586 ( .A(n_466), .B(n_545), .Y(n_586) );
BUFx2_ASAP7_75t_L g718 ( .A(n_466), .Y(n_718) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g487 ( .A(n_467), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g568 ( .A(n_467), .B(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_476), .Y(n_621) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_467), .Y(n_657) );
AND2x2_ASAP7_75t_L g544 ( .A(n_476), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_SL g556 ( .A(n_476), .Y(n_556) );
INVx2_ASAP7_75t_L g567 ( .A(n_476), .Y(n_567) );
BUFx2_ASAP7_75t_L g591 ( .A(n_476), .Y(n_591) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_476), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
AOI332xp33_ASAP7_75t_L g569 ( .A1(n_485), .A2(n_570), .A3(n_574), .B1(n_575), .B2(n_579), .B3(n_582), .C1(n_583), .C2(n_585), .Y(n_569) );
NAND2x1_ASAP7_75t_L g654 ( .A(n_485), .B(n_545), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_485), .B(n_559), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_SL g587 ( .A1(n_486), .A2(n_588), .B(n_591), .C(n_592), .Y(n_587) );
AND2x2_ASAP7_75t_L g726 ( .A(n_486), .B(n_567), .Y(n_726) );
INVx3_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g623 ( .A(n_487), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g628 ( .A(n_487), .B(n_625), .Y(n_628) );
INVx1_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
AND2x2_ASAP7_75t_L g662 ( .A(n_488), .B(n_621), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_488), .B(n_602), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_488), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_488), .B(n_580), .Y(n_688) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g727 ( .A1(n_499), .A2(n_648), .A3(n_655), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
AND2x2_ASAP7_75t_L g531 ( .A(n_500), .B(n_532), .Y(n_531) );
NAND2x1_ASAP7_75t_SL g550 ( .A(n_500), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_500), .Y(n_637) );
AND2x2_ASAP7_75t_L g642 ( .A(n_500), .B(n_553), .Y(n_642) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_501), .A2(n_555), .B(n_557), .C(n_560), .Y(n_554) );
OR2x2_ASAP7_75t_L g571 ( .A(n_501), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
AND2x2_ASAP7_75t_L g590 ( .A(n_501), .B(n_533), .Y(n_590) );
INVx2_ASAP7_75t_L g608 ( .A(n_501), .Y(n_608) );
AND2x2_ASAP7_75t_L g619 ( .A(n_501), .B(n_573), .Y(n_619) );
AND2x2_ASAP7_75t_L g651 ( .A(n_501), .B(n_609), .Y(n_651) );
AND2x2_ASAP7_75t_L g655 ( .A(n_501), .B(n_578), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_501), .B(n_510), .Y(n_660) );
AND2x2_ASAP7_75t_L g694 ( .A(n_501), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_501), .B(n_597), .Y(n_728) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_510), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g636 ( .A(n_510), .Y(n_636) );
AND2x2_ASAP7_75t_L g698 ( .A(n_510), .B(n_619), .Y(n_698) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
OR2x2_ASAP7_75t_L g552 ( .A(n_511), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g562 ( .A(n_511), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g670 ( .A(n_511), .Y(n_670) );
AND2x2_ASAP7_75t_L g687 ( .A(n_511), .B(n_533), .Y(n_687) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g578 ( .A(n_512), .B(n_522), .Y(n_578) );
AND2x2_ASAP7_75t_L g607 ( .A(n_512), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g618 ( .A(n_512), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_512), .B(n_573), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g532 ( .A(n_523), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
AND2x2_ASAP7_75t_L g609 ( .A(n_523), .B(n_573), .Y(n_609) );
INVx1_ASAP7_75t_L g711 ( .A(n_531), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_532), .Y(n_715) );
INVx2_ASAP7_75t_L g573 ( .A(n_533), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_544), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_544), .B(n_649), .Y(n_707) );
OR2x2_ASAP7_75t_L g548 ( .A(n_545), .B(n_546), .Y(n_548) );
INVx1_ASAP7_75t_SL g600 ( .A(n_545), .Y(n_600) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_551), .A2(n_604), .B1(n_606), .B2(n_610), .C(n_611), .Y(n_603) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g631 ( .A(n_552), .B(n_595), .Y(n_631) );
INVx2_ASAP7_75t_L g563 ( .A(n_553), .Y(n_563) );
INVx1_ASAP7_75t_L g589 ( .A(n_553), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_553), .B(n_573), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_553), .B(n_576), .Y(n_683) );
INVx1_ASAP7_75t_L g691 ( .A(n_553), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_555), .B(n_559), .Y(n_605) );
AND2x4_ASAP7_75t_L g580 ( .A(n_556), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g693 ( .A(n_559), .B(n_649), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_562), .B(n_594), .Y(n_593) );
INVxp67_ASAP7_75t_L g701 ( .A(n_563), .Y(n_701) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g601 ( .A(n_567), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g673 ( .A(n_567), .B(n_649), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_567), .B(n_586), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g633 ( .A1(n_568), .A2(n_602), .A3(n_609), .B1(n_634), .B2(n_637), .C1(n_638), .C2(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_568), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g699 ( .A(n_571), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g645 ( .A(n_572), .Y(n_645) );
INVx2_ASAP7_75t_L g576 ( .A(n_573), .Y(n_576) );
INVx1_ASAP7_75t_L g635 ( .A(n_573), .Y(n_635) );
CKINVDCx16_ASAP7_75t_R g582 ( .A(n_574), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g671 ( .A(n_576), .B(n_584), .Y(n_671) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g583 ( .A(n_578), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g626 ( .A(n_578), .B(n_619), .Y(n_626) );
AND2x2_ASAP7_75t_L g630 ( .A(n_578), .B(n_590), .Y(n_630) );
OAI21xp33_ASAP7_75t_SL g640 ( .A1(n_579), .A2(n_641), .B(n_643), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_579), .A2(n_711), .B1(n_712), .B2(n_714), .Y(n_710) );
INVx3_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g585 ( .A(n_580), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_580), .B(n_600), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_582), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g722 ( .A(n_589), .Y(n_722) );
INVx4_ASAP7_75t_L g595 ( .A(n_590), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_590), .B(n_617), .Y(n_665) );
INVx1_ASAP7_75t_SL g677 ( .A(n_591), .Y(n_677) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_595), .B(n_691), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B(n_603), .C(n_620), .Y(n_596) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_598), .A2(n_636), .B1(n_715), .B2(n_717), .C(n_719), .Y(n_716) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_600), .B(n_713), .Y(n_712) );
OAI31xp33_ASAP7_75t_L g692 ( .A1(n_601), .A2(n_678), .A3(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g632 ( .A(n_602), .Y(n_632) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g682 ( .A(n_607), .Y(n_682) );
AND2x2_ASAP7_75t_L g695 ( .A(n_609), .B(n_618), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_615), .Y(n_611) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_619), .B(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_629), .B1(n_631), .B2(n_632), .C(n_633), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_628), .A2(n_697), .B(n_699), .C(n_702), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_631), .B(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g658 ( .A(n_639), .Y(n_658) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_642), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_642), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B(n_652), .C(n_661), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_650), .A2(n_660), .B1(n_724), .B2(n_725), .C(n_727), .Y(n_723) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_656), .B2(n_659), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_SL g724 ( .A(n_663), .Y(n_724) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_696), .C(n_716), .D(n_723), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_672), .B(n_674), .C(n_692), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B(n_680), .C(n_684), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g703 ( .A(n_681), .Y(n_703) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OR2x2_ASAP7_75t_L g714 ( .A(n_682), .B(n_715), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_706), .B2(n_708), .C(n_710), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_713), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_741), .Y(n_745) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
endmodule