module fake_jpeg_25617_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_1),
.B(n_5),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_13),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_23),
.Y(n_44)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_28),
.B1(n_32),
.B2(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_28),
.B1(n_31),
.B2(n_12),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_17),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_14),
.B(n_15),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_61),
.B(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_18),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_60),
.B(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_24),
.B(n_15),
.C(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_55),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_66),
.C(n_57),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_31),
.C(n_7),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_1),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_64),
.Y(n_91)
);

NOR4xp25_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_59),
.C(n_52),
.D(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_11),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_50),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_47),
.B1(n_58),
.B2(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_105),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_80),
.B(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_73),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.C(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_69),
.C(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_94),
.Y(n_106)
);

AO221x1_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_84),
.B1(n_80),
.B2(n_81),
.C(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_83),
.C(n_72),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_112),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_69),
.B1(n_73),
.B2(n_9),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_105),
.B(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_117),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_101),
.B(n_112),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_106),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_111),
.B1(n_99),
.B2(n_114),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_125),
.B1(n_118),
.B2(n_3),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_123),
.B(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_128),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_8),
.C(n_10),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_127),
.C(n_11),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_133),
.B(n_4),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_2),
.B(n_3),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);


endmodule