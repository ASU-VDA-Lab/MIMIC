module real_jpeg_29358_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_9),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_41),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_9),
.B1(n_43),
.B2(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_9),
.B(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_64),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_8),
.A2(n_10),
.B(n_36),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_8),
.A2(n_22),
.B(n_37),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_47),
.Y(n_173)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_10),
.B1(n_48),
.B2(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_9),
.A2(n_43),
.B(n_150),
.C(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_118),
.CON(n_12),
.SN(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_99),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_15),
.B(n_99),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_79),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_68),
.B2(n_69),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_20),
.A2(n_32),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_20),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_21),
.B(n_24),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_21),
.A2(n_29),
.B1(n_86),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_27),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_29),
.A2(n_83),
.B(n_112),
.Y(n_140)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_29),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_32),
.A2(n_103),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_32),
.A2(n_103),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_32),
.B(n_111),
.C(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_32),
.B(n_156),
.C(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_33),
.B(n_39),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_36),
.A2(n_38),
.B(n_43),
.C(n_170),
.Y(n_169)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_39),
.B(n_43),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_59),
.B(n_62),
.C(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_43),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_45),
.B(n_96),
.C(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_45),
.A2(n_66),
.B1(n_126),
.B2(n_127),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_45),
.A2(n_66),
.B1(n_87),
.B2(n_88),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_51),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_46),
.A2(n_49),
.B1(n_94),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_107),
.C(n_113),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_55),
.A2(n_67),
.B1(n_113),
.B2(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_88),
.C(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_77),
.B(n_85),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.C(n_95),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_87),
.B1(n_88),
.B2(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_87),
.A2(n_88),
.B1(n_169),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_88),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_96),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_100),
.B(n_102),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_105),
.A2(n_106),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_111),
.A2(n_138),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_187),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_114),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_140),
.C(n_141),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_143),
.B(n_203),
.C(n_208),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_133),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_120),
.B(n_133),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_124),
.C(n_131),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_134),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_139),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_140),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_202),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_197),
.B(n_201),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_165),
.B(n_196),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_147),
.B(n_155),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_154),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_191),
.B(n_195),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_176),
.B(n_190),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B(n_189),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_188),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);


endmodule