module fake_ariane_2048_n_1724 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1724);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1724;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_44),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_21),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_40),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_29),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_85),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_80),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_81),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_101),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_28),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_61),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_57),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_28),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_47),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_2),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_87),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_44),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_4),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_1),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_13),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_6),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_24),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_46),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_20),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_70),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_15),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_12),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_74),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_53),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_113),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_48),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_86),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_112),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_127),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_141),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_54),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_51),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_51),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_110),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_38),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_45),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_43),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_18),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_107),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_124),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_103),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_137),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_84),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_36),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_24),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_92),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_41),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_116),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_23),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_114),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_72),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_122),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_96),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_42),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_125),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_105),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_97),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_66),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_17),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_88),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_18),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_8),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_71),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_35),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_78),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_32),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_8),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_47),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_52),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_33),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_150),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_98),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_43),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_34),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_152),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_169),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_161),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_174),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_161),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_291),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_169),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_162),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_165),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_186),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_162),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_163),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_233),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_235),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_168),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_187),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_175),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_175),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_178),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_221),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_209),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_221),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_178),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_269),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_189),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_194),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_157),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_157),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_269),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_183),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_183),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_204),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_184),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_216),
.B(n_0),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_198),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_151),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_216),
.B(n_2),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_167),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_157),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_226),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_198),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_176),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_177),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_180),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_208),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_208),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_191),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_215),
.B(n_3),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_215),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_219),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_176),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_219),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_192),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_243),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_195),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_220),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_186),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_220),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_225),
.B(n_4),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_278),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_196),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_201),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_176),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_158),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_156),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_309),
.B(n_200),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_245),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_320),
.A2(n_193),
.B1(n_272),
.B2(n_292),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_302),
.B(n_252),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_304),
.B(n_203),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_304),
.B(n_252),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_339),
.B(n_164),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_342),
.B(n_228),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_307),
.B(n_261),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_310),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_312),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_316),
.A2(n_265),
.B(n_261),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_329),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_276),
.B(n_228),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_350),
.B(n_265),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_335),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

AND3x2_ASAP7_75t_L g423 ( 
.A(n_306),
.B(n_237),
.C(n_203),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_156),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_203),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_346),
.B(n_156),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_346),
.B(n_271),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_351),
.B(n_271),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_348),
.B(n_237),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_341),
.B(n_343),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_356),
.B(n_230),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_309),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_393),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_388),
.B(n_363),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_440),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_363),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_332),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_276),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_344),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_376),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_418),
.B(n_349),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_418),
.B(n_353),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_359),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_395),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_318),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_385),
.B(n_361),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_377),
.B(n_357),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_R g468 ( 
.A(n_387),
.B(n_301),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_276),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_438),
.B(n_371),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_374),
.A2(n_354),
.B1(n_193),
.B2(n_272),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_358),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_358),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_377),
.B(n_362),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_440),
.B(n_368),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_374),
.B(n_370),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_392),
.B(n_373),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_277),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_377),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_381),
.B(n_362),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_381),
.B(n_364),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_419),
.B(n_364),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g499 ( 
.A1(n_409),
.A2(n_366),
.B(n_283),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_365),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_396),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_396),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_396),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

CKINVDCx6p67_ASAP7_75t_R g512 ( 
.A(n_404),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_365),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_437),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_425),
.B(n_164),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_419),
.B(n_369),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_419),
.B(n_369),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_391),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_379),
.A2(n_325),
.B1(n_299),
.B2(n_213),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_379),
.B(n_213),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_425),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_402),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_381),
.B(n_155),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

INVx8_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_425),
.A2(n_237),
.B1(n_155),
.B2(n_297),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_411),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_424),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_392),
.B(n_372),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_389),
.B(n_283),
.C(n_277),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_384),
.B(n_303),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_394),
.B(n_398),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_411),
.A2(n_207),
.B1(n_240),
.B2(n_236),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_424),
.B(n_200),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_424),
.B(n_287),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_416),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_425),
.A2(n_206),
.B1(n_223),
.B2(n_218),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_287),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_384),
.B(n_210),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_381),
.B(n_181),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_394),
.B(n_308),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_398),
.B(n_313),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_416),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_395),
.B(n_305),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_425),
.B(n_164),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_402),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_378),
.A2(n_275),
.B1(n_242),
.B2(n_297),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_430),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_434),
.B(n_275),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_432),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_412),
.B(n_314),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_381),
.B(n_181),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_432),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_432),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_399),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_412),
.B(n_211),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_434),
.B(n_153),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_432),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_414),
.B(n_224),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_442),
.A2(n_223),
.B1(n_242),
.B2(n_249),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_381),
.B(n_185),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_439),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_426),
.B(n_185),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_404),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_462),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_446),
.B(n_434),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_R g595 ( 
.A(n_468),
.B(n_330),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_462),
.Y(n_596)
);

AO22x2_ASAP7_75t_L g597 ( 
.A1(n_448),
.A2(n_188),
.B1(n_202),
.B2(n_206),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_444),
.B(n_470),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_L g599 ( 
.A(n_444),
.B(n_439),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_434),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_460),
.A2(n_442),
.B1(n_425),
.B2(n_429),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_450),
.A2(n_434),
.B(n_406),
.C(n_422),
.Y(n_603)
);

OAI221xp5_ASAP7_75t_L g604 ( 
.A1(n_473),
.A2(n_202),
.B1(n_188),
.B2(n_212),
.C(n_214),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_474),
.B(n_389),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_489),
.B(n_378),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_576),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_466),
.B(n_389),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_474),
.B(n_401),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_451),
.A2(n_402),
.B1(n_442),
.B2(n_429),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_458),
.B(n_401),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_451),
.A2(n_402),
.B1(n_442),
.B2(n_429),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_536),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_476),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_474),
.B(n_401),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_405),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_536),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_480),
.B(n_405),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_455),
.A2(n_442),
.B1(n_425),
.B2(n_429),
.Y(n_620)
);

OAI221xp5_ASAP7_75t_L g621 ( 
.A1(n_473),
.A2(n_238),
.B1(n_292),
.B2(n_256),
.C(n_255),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_480),
.A2(n_442),
.B1(n_429),
.B2(n_417),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_380),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_453),
.B(n_439),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_451),
.A2(n_402),
.B1(n_429),
.B2(n_442),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_540),
.Y(n_626)
);

BUFx5_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_464),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_423),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_528),
.A2(n_390),
.B1(n_431),
.B2(n_380),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_480),
.B(n_406),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_447),
.B(n_541),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g633 ( 
.A(n_443),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_508),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_447),
.B(n_406),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_540),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_453),
.B(n_415),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_461),
.B(n_214),
.C(n_212),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_518),
.B(n_402),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_540),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_464),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_578),
.B(n_415),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_415),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_465),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_511),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_487),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_494),
.B(n_422),
.Y(n_647)
);

AND2x2_ASAP7_75t_SL g648 ( 
.A(n_518),
.B(n_383),
.Y(n_648)
);

BUFx6f_ASAP7_75t_SL g649 ( 
.A(n_528),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_490),
.B(n_383),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_519),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_453),
.B(n_520),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_453),
.B(n_520),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_494),
.B(n_422),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_520),
.B(n_529),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_488),
.B(n_417),
.Y(n_656)
);

BUFx5_ASAP7_75t_L g657 ( 
.A(n_484),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_465),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_496),
.B(n_420),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_524),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_539),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_524),
.Y(n_663)
);

AO22x1_ASAP7_75t_L g664 ( 
.A1(n_461),
.A2(n_442),
.B1(n_429),
.B2(n_426),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_447),
.B(n_420),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_447),
.B(n_421),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_539),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_471),
.B(n_421),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_520),
.B(n_427),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_471),
.B(n_427),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_544),
.B(n_441),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_452),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_467),
.B(n_441),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_445),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_484),
.B(n_423),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_547),
.B(n_449),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_443),
.B(n_390),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_556),
.B(n_431),
.Y(n_678)
);

BUFx6f_ASAP7_75t_SL g679 ( 
.A(n_528),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_557),
.B(n_433),
.C(n_400),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_571),
.B(n_433),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_452),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_454),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_449),
.B(n_397),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_449),
.B(n_397),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_528),
.B(n_336),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_492),
.B(n_397),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_456),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_516),
.B(n_397),
.Y(n_689)
);

BUFx12f_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_492),
.B(n_400),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_492),
.B(n_400),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_487),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_451),
.A2(n_442),
.B1(n_429),
.B2(n_426),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_529),
.B(n_400),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_456),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_498),
.A2(n_436),
.B(n_435),
.C(n_403),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_454),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_500),
.A2(n_436),
.B(n_435),
.C(n_403),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_457),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_483),
.B(n_403),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_515),
.B(n_403),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_472),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_522),
.B(n_408),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_563),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_516),
.B(n_426),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_472),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_457),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_561),
.A2(n_442),
.B1(n_429),
.B2(n_426),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_546),
.B(n_413),
.C(n_408),
.Y(n_710)
);

CKINVDCx14_ASAP7_75t_R g711 ( 
.A(n_512),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_529),
.B(n_408),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_561),
.A2(n_429),
.B1(n_426),
.B2(n_435),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_475),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_475),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_563),
.B(n_386),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_529),
.B(n_408),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_523),
.B(n_413),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_463),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_548),
.A2(n_436),
.B(n_435),
.C(n_428),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_477),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_560),
.B(n_444),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_477),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_463),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_451),
.A2(n_429),
.B1(n_436),
.B2(n_428),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_531),
.B(n_413),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_531),
.B(n_413),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_555),
.B(n_428),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_554),
.B(n_428),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_481),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_555),
.B(n_386),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_525),
.A2(n_217),
.B1(n_218),
.B2(n_238),
.C(n_241),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_528),
.A2(n_256),
.B1(n_241),
.B2(n_249),
.Y(n_733)
);

AO22x1_ASAP7_75t_L g734 ( 
.A1(n_491),
.A2(n_253),
.B1(n_262),
.B2(n_264),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_478),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_586),
.B(n_386),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_478),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_579),
.A2(n_409),
.B(n_386),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_479),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_591),
.B(n_409),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_586),
.B(n_386),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_487),
.B(n_229),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_481),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_479),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_572),
.B(n_217),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_560),
.B(n_154),
.Y(n_746)
);

INVxp33_ASAP7_75t_L g747 ( 
.A(n_543),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_590),
.B(n_251),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_560),
.B(n_159),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_590),
.B(n_251),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_572),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_491),
.A2(n_171),
.B1(n_170),
.B2(n_166),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_487),
.B(n_232),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_572),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_572),
.B(n_244),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_560),
.B(n_160),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_527),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_444),
.B(n_172),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_676),
.A2(n_691),
.B(n_684),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_662),
.B(n_525),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_678),
.B(n_681),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_662),
.B(n_345),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_632),
.B(n_590),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_668),
.B(n_590),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_630),
.A2(n_650),
.B1(n_606),
.B2(n_592),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_637),
.A2(n_562),
.B(n_530),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_668),
.B(n_491),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_665),
.B(n_491),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_672),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_682),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_738),
.A2(n_562),
.B(n_530),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_665),
.B(n_491),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_637),
.A2(n_486),
.B(n_485),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_642),
.B(n_534),
.Y(n_775)
);

O2A1O1Ixp5_ASAP7_75t_L g776 ( 
.A1(n_608),
.A2(n_567),
.B(n_552),
.C(n_549),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_688),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_754),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_623),
.B(n_542),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_754),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_674),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_594),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_593),
.A2(n_486),
.B(n_485),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_594),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_669),
.A2(n_502),
.B(n_495),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_633),
.B(n_504),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_594),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_666),
.A2(n_542),
.B(n_259),
.C(n_267),
.Y(n_788)
);

INVx11_ASAP7_75t_L g789 ( 
.A(n_690),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_596),
.B(n_677),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_594),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_630),
.B(n_444),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_666),
.B(n_491),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_669),
.A2(n_502),
.B(n_495),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_670),
.B(n_491),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_696),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_701),
.A2(n_505),
.B(n_497),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_605),
.A2(n_255),
.B(n_259),
.C(n_267),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_595),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_667),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_700),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_611),
.B(n_451),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_628),
.B(n_360),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_611),
.B(n_451),
.Y(n_804)
);

AOI21xp33_ASAP7_75t_L g805 ( 
.A1(n_607),
.A2(n_565),
.B(n_550),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_617),
.B(n_469),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_617),
.A2(n_673),
.B(n_656),
.C(n_616),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_643),
.A2(n_583),
.B1(n_534),
.B2(n_538),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_624),
.A2(n_687),
.B(n_685),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_624),
.A2(n_505),
.B(n_497),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_636),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_656),
.B(n_469),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_685),
.A2(n_501),
.B(n_482),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_708),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_595),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_751),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_671),
.B(n_469),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_641),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_673),
.B(n_609),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_687),
.A2(n_501),
.B(n_482),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_619),
.A2(n_286),
.B(n_588),
.C(n_587),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_692),
.A2(n_506),
.B(n_503),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_719),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_631),
.A2(n_286),
.B(n_588),
.C(n_587),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_733),
.A2(n_565),
.B1(n_469),
.B2(n_534),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_742),
.B(n_469),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_695),
.A2(n_506),
.B(n_503),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_629),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_648),
.B(n_470),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_644),
.B(n_504),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_692),
.A2(n_509),
.B(n_507),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_742),
.B(n_469),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_695),
.A2(n_509),
.B(n_507),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_711),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_712),
.A2(n_514),
.B(n_510),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_724),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_753),
.B(n_565),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_648),
.A2(n_600),
.B1(n_654),
.B2(n_647),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_753),
.B(n_565),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_735),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_L g841 ( 
.A1(n_758),
.A2(n_504),
.B(n_513),
.C(n_526),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_712),
.A2(n_568),
.B(n_558),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_717),
.A2(n_551),
.B(n_514),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_758),
.A2(n_513),
.B(n_526),
.C(n_549),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_659),
.B(n_470),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_639),
.B(n_470),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_636),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_639),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_627),
.B(n_534),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_658),
.B(n_513),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_627),
.B(n_534),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_733),
.A2(n_559),
.B1(n_549),
.B2(n_526),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_733),
.A2(n_517),
.B1(n_535),
.B2(n_584),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_717),
.A2(n_517),
.B(n_535),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_737),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_601),
.B(n_470),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_706),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_629),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_716),
.B(n_545),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_680),
.B(n_493),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_747),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_702),
.A2(n_558),
.B(n_545),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_755),
.B(n_493),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_726),
.A2(n_551),
.B1(n_564),
.B2(n_573),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_683),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_739),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_622),
.B(n_493),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_698),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_703),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_704),
.A2(n_573),
.B(n_564),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_707),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_638),
.B(n_367),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_746),
.A2(n_574),
.B(n_575),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_718),
.A2(n_574),
.B(n_575),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_722),
.A2(n_577),
.B(n_585),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_714),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_706),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_722),
.A2(n_577),
.B(n_585),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_598),
.A2(n_589),
.B(n_527),
.Y(n_879)
);

AO21x1_ASAP7_75t_L g880 ( 
.A1(n_720),
.A2(n_589),
.B(n_532),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_649),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_744),
.Y(n_882)
);

CKINVDCx14_ASAP7_75t_R g883 ( 
.A(n_675),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_635),
.A2(n_537),
.B(n_580),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_604),
.A2(n_580),
.B(n_570),
.C(n_532),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_646),
.B(n_493),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_746),
.A2(n_537),
.B(n_570),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_731),
.A2(n_736),
.B(n_741),
.C(n_728),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_755),
.B(n_493),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_749),
.A2(n_553),
.B(n_533),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_614),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_686),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_740),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_706),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_715),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_749),
.A2(n_553),
.B(n_533),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_729),
.B(n_521),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_756),
.A2(n_499),
.B(n_521),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_756),
.A2(n_499),
.B(n_521),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_652),
.A2(n_499),
.B(n_521),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_697),
.A2(n_581),
.B(n_521),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_627),
.B(n_569),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_699),
.A2(n_581),
.B(n_230),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_729),
.B(n_745),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_646),
.B(n_581),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_721),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_748),
.B(n_581),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_634),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_652),
.A2(n_581),
.B(n_569),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_602),
.B(n_569),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_258),
.B1(n_298),
.B2(n_296),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_750),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_723),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_693),
.B(n_569),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_706),
.A2(n_569),
.B1(n_295),
.B2(n_279),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_613),
.B(n_569),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_618),
.B(n_281),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_653),
.A2(n_294),
.B(n_293),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_740),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_603),
.A2(n_290),
.B(n_282),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_653),
.A2(n_285),
.B(n_173),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_740),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_597),
.B(n_730),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_655),
.A2(n_239),
.B(n_280),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_655),
.A2(n_234),
.B(n_274),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_599),
.A2(n_231),
.B(n_273),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_706),
.B(n_284),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_743),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_757),
.A2(n_270),
.B(n_268),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_693),
.B(n_263),
.Y(n_930)
);

AOI33xp33_ASAP7_75t_L g931 ( 
.A1(n_626),
.A2(n_7),
.A3(n_15),
.B1(n_20),
.B2(n_21),
.B3(n_22),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_640),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_645),
.A2(n_260),
.B(n_257),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_710),
.A2(n_660),
.B(n_663),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_732),
.A2(n_230),
.B(n_250),
.Y(n_935)
);

AND2x2_ASAP7_75t_SL g936 ( 
.A(n_610),
.B(n_164),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_651),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_661),
.A2(n_248),
.B(n_247),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_627),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_689),
.A2(n_246),
.B(n_227),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_664),
.A2(n_222),
.B(n_205),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_762),
.B(n_621),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_781),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_828),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_807),
.A2(n_615),
.B(n_725),
.C(n_612),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_764),
.B(n_597),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_790),
.B(n_597),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_765),
.B(n_694),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_807),
.A2(n_725),
.B(n_612),
.C(n_625),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_789),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_SL g951 ( 
.A(n_834),
.B(n_179),
.C(n_182),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_803),
.A2(n_679),
.B1(n_649),
.B2(n_734),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_761),
.A2(n_709),
.B(n_713),
.C(n_620),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_760),
.B(n_679),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_799),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_761),
.A2(n_752),
.B(n_610),
.C(n_625),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_819),
.A2(n_772),
.B(n_775),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_920),
.B(n_694),
.C(n_199),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_790),
.B(n_657),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_809),
.A2(n_657),
.B(n_627),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_SL g961 ( 
.A1(n_859),
.A2(n_7),
.B(n_22),
.C(n_23),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_936),
.A2(n_657),
.B1(n_627),
.B2(n_197),
.Y(n_962)
);

AO32x2_ASAP7_75t_L g963 ( 
.A1(n_838),
.A2(n_657),
.A3(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_759),
.A2(n_657),
.B(n_190),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_770),
.B(n_25),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_849),
.A2(n_25),
.B(n_27),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_788),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_788),
.A2(n_911),
.B(n_763),
.C(n_778),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_903),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_800),
.B(n_818),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_851),
.A2(n_36),
.B(n_37),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_828),
.B(n_37),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_38),
.B(n_39),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_778),
.B(n_41),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_936),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_859),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_792),
.A2(n_55),
.B(n_56),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_898),
.A2(n_90),
.B(n_142),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_861),
.B(n_57),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_888),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_821),
.A2(n_59),
.B(n_64),
.C(n_65),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_912),
.B(n_67),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_865),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_780),
.B(n_69),
.Y(n_984)
);

AND2x4_ASAP7_75t_SL g985 ( 
.A(n_815),
.B(n_82),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_816),
.B(n_89),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_868),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_SL g988 ( 
.A(n_917),
.B(n_95),
.C(n_100),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_763),
.A2(n_102),
.B(n_118),
.C(n_119),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_L g990 ( 
.A1(n_901),
.A2(n_120),
.B(n_121),
.C(n_135),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_931),
.B(n_136),
.C(n_144),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_858),
.B(n_857),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_892),
.B(n_872),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_816),
.A2(n_779),
.B1(n_919),
.B2(n_786),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_857),
.B(n_877),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_869),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_904),
.B(n_858),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_900),
.A2(n_890),
.B(n_887),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_881),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_824),
.B(n_798),
.C(n_889),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_786),
.B(n_830),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_883),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_857),
.B(n_877),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_824),
.A2(n_863),
.B(n_767),
.C(n_906),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_845),
.A2(n_773),
.B(n_768),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_882),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_883),
.B(n_923),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_937),
.B(n_782),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_850),
.A2(n_917),
.B(n_871),
.C(n_913),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_793),
.A2(n_817),
.B(n_783),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_847),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_797),
.A2(n_832),
.B(n_826),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_877),
.B(n_894),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_847),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_876),
.A2(n_895),
.B1(n_928),
.B2(n_808),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_769),
.Y(n_1017)
);

BUFx8_ASAP7_75t_L g1018 ( 
.A(n_877),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_931),
.B(n_937),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_795),
.A2(n_812),
.B(n_804),
.C(n_802),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_805),
.B(n_837),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_856),
.A2(n_874),
.B(n_870),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_811),
.A2(n_806),
.B1(n_825),
.B2(n_839),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_811),
.B(n_825),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_893),
.A2(n_922),
.B1(n_907),
.B2(n_864),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_771),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_856),
.A2(n_862),
.B(n_897),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_777),
.Y(n_1028)
);

AOI22x1_ASAP7_75t_L g1029 ( 
.A1(n_813),
.A2(n_822),
.B1(n_820),
.B2(n_831),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_852),
.B(n_932),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_922),
.B(n_935),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_847),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_885),
.A2(n_829),
.B(n_934),
.C(n_853),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_927),
.A2(n_860),
.B(n_930),
.C(n_867),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_896),
.A2(n_785),
.B(n_794),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_899),
.A2(n_879),
.B(n_873),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_847),
.B(n_894),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_796),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_782),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_774),
.A2(n_810),
.B(n_878),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_894),
.A2(n_932),
.B1(n_848),
.B2(n_915),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_801),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_894),
.B(n_848),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_766),
.A2(n_776),
.B(n_841),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_867),
.A2(n_910),
.B(n_916),
.C(n_844),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_814),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_910),
.A2(n_916),
.B(n_846),
.C(n_939),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_902),
.B(n_932),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_836),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_932),
.B(n_848),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_875),
.A2(n_884),
.B(n_846),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_840),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_855),
.B(n_908),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_782),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_930),
.A2(n_886),
.B(n_905),
.C(n_827),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_866),
.B(n_891),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_782),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_791),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_902),
.B(n_939),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_784),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_787),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_787),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_791),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_933),
.A2(n_940),
.B1(n_914),
.B2(n_921),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_833),
.A2(n_835),
.B(n_842),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_905),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_918),
.B(n_925),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_843),
.A2(n_854),
.B(n_880),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_924),
.A2(n_914),
.B1(n_938),
.B2(n_929),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_941),
.B(n_926),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_909),
.B(n_650),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_SL g1073 ( 
.A1(n_936),
.A2(n_648),
.B(n_764),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_L g1074 ( 
.A(n_819),
.B(n_807),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_823),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_762),
.B(n_591),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_SL g1077 ( 
.A(n_834),
.B(n_488),
.C(n_559),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_823),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_803),
.B(n_461),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_L g1080 ( 
.A(n_761),
.B(n_461),
.C(n_632),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_807),
.A2(n_466),
.B(n_460),
.C(n_765),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_1081),
.B(n_1074),
.C(n_975),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_943),
.Y(n_1083)
);

BUFx10_ASAP7_75t_L g1084 ( 
.A(n_950),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1079),
.B(n_970),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_942),
.B(n_1008),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_957),
.A2(n_1060),
.B(n_960),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_L g1088 ( 
.A(n_980),
.B(n_977),
.C(n_973),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_957),
.A2(n_960),
.B(n_1048),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1073),
.A2(n_948),
.B1(n_1019),
.B2(n_976),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1005),
.A2(n_1035),
.B(n_1022),
.Y(n_1092)
);

AO21x1_ASAP7_75t_L g1093 ( 
.A1(n_980),
.A2(n_977),
.B(n_973),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1076),
.B(n_954),
.Y(n_1094)
);

AOI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_968),
.A2(n_949),
.B(n_1000),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_994),
.B(n_955),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1005),
.A2(n_1035),
.B(n_964),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_961),
.A2(n_965),
.B(n_972),
.C(n_1010),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1051),
.A2(n_998),
.B(n_1040),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1002),
.Y(n_1100)
);

AND2x6_ASAP7_75t_SL g1101 ( 
.A(n_974),
.B(n_947),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_964),
.A2(n_1013),
.B(n_1011),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_997),
.B(n_983),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1020),
.A2(n_953),
.B(n_1004),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_956),
.A2(n_945),
.B(n_958),
.C(n_1000),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1047),
.A2(n_1045),
.B(n_1040),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_993),
.B(n_979),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_987),
.B(n_996),
.Y(n_1108)
);

AOI221x1_ASAP7_75t_L g1109 ( 
.A1(n_966),
.A2(n_971),
.B1(n_991),
.B2(n_1069),
.C(n_1025),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_999),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1027),
.A2(n_1066),
.B(n_1029),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1034),
.A2(n_1030),
.B(n_981),
.C(n_971),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_967),
.A2(n_981),
.B(n_1001),
.C(n_966),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_1016),
.A2(n_1034),
.B(n_962),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_944),
.B(n_1012),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1077),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1038),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_959),
.A2(n_1055),
.B(n_984),
.C(n_986),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1046),
.B(n_946),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1021),
.B(n_1050),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1072),
.A2(n_1069),
.B(n_1027),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_SL g1123 ( 
.A1(n_1055),
.A2(n_1057),
.B(n_1068),
.C(n_1033),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1004),
.A2(n_969),
.B(n_988),
.C(n_989),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1023),
.A2(n_1070),
.A3(n_1041),
.B(n_1024),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1044),
.A2(n_990),
.B(n_978),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1015),
.B(n_1018),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1058),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1065),
.A2(n_995),
.B(n_1003),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1043),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1017),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1009),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1042),
.B(n_1049),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_1014),
.A2(n_1037),
.B(n_982),
.C(n_1061),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_992),
.B1(n_1062),
.B2(n_1063),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1006),
.A2(n_1056),
.B(n_1053),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1006),
.A2(n_985),
.B(n_1064),
.C(n_951),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1007),
.A2(n_1078),
.B(n_1075),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_978),
.A2(n_992),
.B(n_1059),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1067),
.A2(n_1059),
.B(n_1032),
.C(n_1052),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_963),
.A2(n_1067),
.A3(n_1043),
.B(n_1058),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1067),
.B(n_1039),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1058),
.A2(n_1039),
.B(n_1054),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_SL g1144 ( 
.A1(n_963),
.A2(n_1039),
.B(n_1054),
.C(n_1058),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1054),
.B(n_963),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_998),
.A2(n_1035),
.B(n_1036),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_942),
.B(n_760),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1002),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_950),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_998),
.A2(n_1035),
.B(n_1036),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_944),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_950),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_SL g1154 ( 
.A(n_1080),
.B(n_395),
.C(n_461),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_998),
.A2(n_1035),
.B(n_1036),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1081),
.A2(n_1073),
.B(n_466),
.C(n_460),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_943),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_942),
.B(n_760),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1081),
.A2(n_632),
.B(n_459),
.C(n_458),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1073),
.B(n_936),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1073),
.A2(n_374),
.B1(n_686),
.B2(n_313),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_998),
.A2(n_1035),
.B(n_1036),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_943),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1081),
.A2(n_807),
.B(n_1005),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1081),
.A2(n_1073),
.B(n_466),
.C(n_460),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_944),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_944),
.B(n_858),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_943),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1081),
.A2(n_1073),
.B(n_466),
.C(n_460),
.Y(n_1176)
);

AO32x2_ASAP7_75t_L g1177 ( 
.A1(n_1025),
.A2(n_1023),
.A3(n_1016),
.B1(n_976),
.B2(n_379),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_944),
.B(n_828),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1079),
.B(n_592),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_950),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1081),
.A2(n_1073),
.B(n_466),
.C(n_460),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_943),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1074),
.B(n_807),
.Y(n_1185)
);

AO32x2_ASAP7_75t_L g1186 ( 
.A1(n_1025),
.A2(n_1023),
.A3(n_1016),
.B1(n_976),
.B2(n_379),
.Y(n_1186)
);

NOR4xp25_ASAP7_75t_L g1187 ( 
.A(n_1081),
.B(n_980),
.C(n_975),
.D(n_967),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1081),
.A2(n_807),
.B(n_819),
.C(n_632),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1080),
.B(n_461),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_944),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_944),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_970),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1196)
);

OAI22x1_ASAP7_75t_L g1197 ( 
.A1(n_994),
.A2(n_525),
.B1(n_473),
.B2(n_952),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1081),
.A2(n_632),
.B(n_459),
.C(n_458),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1081),
.A2(n_807),
.B(n_1005),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_L g1201 ( 
.A(n_1058),
.B(n_1006),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1081),
.A2(n_807),
.B(n_819),
.C(n_632),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1081),
.A2(n_807),
.B(n_819),
.C(n_632),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_955),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1002),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1073),
.B(n_936),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_943),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_944),
.B(n_828),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_943),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1081),
.A2(n_807),
.B(n_819),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_942),
.A2(n_936),
.B1(n_374),
.B2(n_528),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1071),
.A2(n_903),
.A3(n_901),
.B(n_880),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_943),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1081),
.A2(n_1074),
.B(n_957),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1036),
.A2(n_1022),
.B(n_1051),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_943),
.Y(n_1220)
);

CKINVDCx11_ASAP7_75t_R g1221 ( 
.A(n_1149),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1132),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1084),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1108),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1181),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1215),
.A2(n_1167),
.B1(n_1197),
.B2(n_1147),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1083),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1121),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1084),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1152),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1117),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1085),
.B(n_1161),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_1086),
.B2(n_1082),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_1082),
.B2(n_1091),
.Y(n_1234)
);

CKINVDCx6p67_ASAP7_75t_R g1235 ( 
.A(n_1110),
.Y(n_1235)
);

BUFx8_ASAP7_75t_L g1236 ( 
.A(n_1148),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1204),
.Y(n_1237)
);

CKINVDCx11_ASAP7_75t_R g1238 ( 
.A(n_1205),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1195),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1154),
.A2(n_1096),
.B1(n_1091),
.B2(n_1179),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1101),
.Y(n_1241)
);

NOR2x1_ASAP7_75t_L g1242 ( 
.A(n_1191),
.B(n_1137),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1127),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1094),
.B(n_1107),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1159),
.A2(n_1171),
.B1(n_1182),
.B2(n_1176),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1128),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_1088),
.B1(n_1185),
.B2(n_1104),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1151),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1095),
.A2(n_1088),
.B1(n_1185),
.B2(n_1104),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1177),
.A2(n_1186),
.B1(n_1145),
.B2(n_1170),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1151),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1160),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1177),
.A2(n_1186),
.B1(n_1170),
.B2(n_1200),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1169),
.B(n_1175),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1177),
.A2(n_1186),
.B1(n_1200),
.B2(n_1121),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1093),
.A2(n_1115),
.B1(n_1103),
.B2(n_1210),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1184),
.A2(n_1208),
.B1(n_1217),
.B2(n_1220),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1213),
.A2(n_1112),
.B1(n_1165),
.B2(n_1199),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1118),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1120),
.B(n_1114),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1100),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1131),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1116),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1133),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1151),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1173),
.A2(n_1101),
.B1(n_1106),
.B2(n_1135),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1113),
.A2(n_1105),
.B1(n_1098),
.B2(n_1218),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1172),
.B(n_1192),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1172),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1138),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1153),
.A2(n_1214),
.B1(n_1190),
.B2(n_1163),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1172),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1155),
.A2(n_1180),
.B1(n_1138),
.B2(n_1187),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1128),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1109),
.A2(n_1130),
.B1(n_1192),
.B2(n_1193),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1124),
.A2(n_1090),
.B1(n_1178),
.B2(n_1209),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1130),
.A2(n_1144),
.B1(n_1141),
.B2(n_1192),
.Y(n_1277)
);

BUFx8_ASAP7_75t_L g1278 ( 
.A(n_1193),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1193),
.A2(n_1142),
.B1(n_1202),
.B2(n_1203),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1136),
.A2(n_1126),
.B1(n_1129),
.B2(n_1139),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1136),
.A2(n_1097),
.B1(n_1189),
.B2(n_1125),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1087),
.A2(n_1140),
.B1(n_1102),
.B2(n_1092),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1201),
.B(n_1123),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1201),
.B(n_1125),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1125),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1134),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1146),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1146),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1111),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1119),
.A2(n_1122),
.B1(n_1157),
.B2(n_1168),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1150),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1150),
.A2(n_1168),
.B1(n_1157),
.B2(n_1099),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1158),
.A2(n_1194),
.B1(n_1216),
.B2(n_1162),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1158),
.A2(n_1194),
.B1(n_1216),
.B2(n_1162),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1162),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1164),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1164),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1219),
.A2(n_1089),
.B1(n_1156),
.B2(n_1212),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1164),
.B(n_1216),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1183),
.A2(n_1194),
.B1(n_1198),
.B2(n_1174),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1183),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1198),
.A2(n_1188),
.B1(n_1196),
.B2(n_1206),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1198),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1211),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1215),
.A2(n_528),
.B1(n_1167),
.B2(n_733),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1215),
.A2(n_528),
.B1(n_1167),
.B2(n_733),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1215),
.A2(n_528),
.B1(n_1167),
.B2(n_733),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1149),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1108),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1195),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1195),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1195),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1181),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1108),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1149),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1132),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1149),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1148),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1195),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1215),
.A2(n_528),
.B1(n_1167),
.B2(n_733),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1195),
.Y(n_1323)
);

BUFx8_ASAP7_75t_SL g1324 ( 
.A(n_1149),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1215),
.A2(n_528),
.B1(n_1167),
.B2(n_733),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_374),
.B2(n_686),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1108),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1108),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1181),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1108),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1121),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1181),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1108),
.Y(n_1333)
);

INVx6_ASAP7_75t_L g1334 ( 
.A(n_1084),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_SL g1335 ( 
.A(n_1149),
.Y(n_1335)
);

INVx11_ASAP7_75t_L g1336 ( 
.A(n_1149),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_374),
.B2(n_686),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_1091),
.B2(n_473),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1181),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1084),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1147),
.B(n_1161),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1084),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1108),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1250),
.B(n_1253),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1319),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1297),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1303),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1282),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1282),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1285),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1286),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1270),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1254),
.B(n_1224),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1324),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1301),
.Y(n_1355)
);

AOI211xp5_ASAP7_75t_L g1356 ( 
.A1(n_1338),
.A2(n_1267),
.B(n_1258),
.C(n_1240),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1298),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1288),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1283),
.A2(n_1293),
.B(n_1271),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1289),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1305),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1245),
.A2(n_1295),
.A3(n_1302),
.B(n_1287),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1228),
.B(n_1331),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_1221),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1311),
.B(n_1316),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1227),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1252),
.Y(n_1368)
);

AO21x1_ASAP7_75t_L g1369 ( 
.A1(n_1338),
.A2(n_1275),
.B(n_1296),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1293),
.A2(n_1271),
.B(n_1300),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1259),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1275),
.A2(n_1304),
.B(n_1306),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1299),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1221),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1290),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1294),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1294),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1247),
.A2(n_1249),
.B(n_1234),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1262),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1314),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1326),
.A2(n_1337),
.B1(n_1308),
.B2(n_1307),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1290),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1222),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1321),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1239),
.Y(n_1385)
);

INVx3_ASAP7_75t_SL g1386 ( 
.A(n_1334),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1312),
.B(n_1313),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1330),
.B(n_1333),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1292),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1222),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1318),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1255),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1323),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1244),
.B(n_1343),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1284),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1264),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1341),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1318),
.Y(n_1398)
);

AOI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1276),
.A2(n_1242),
.B(n_1268),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1260),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1257),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1234),
.A2(n_1233),
.B(n_1309),
.C(n_1307),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1256),
.A2(n_1273),
.B(n_1249),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1246),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1247),
.B(n_1256),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1246),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1273),
.A2(n_1266),
.B(n_1274),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1257),
.B(n_1232),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1263),
.A2(n_1291),
.B(n_1243),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1233),
.B(n_1266),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1226),
.A2(n_1281),
.B(n_1304),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1248),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1308),
.A2(n_1325),
.B(n_1322),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1277),
.A2(n_1280),
.B(n_1226),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1279),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1251),
.B(n_1265),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1241),
.B(n_1237),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1229),
.A2(n_1342),
.B(n_1340),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1310),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1278),
.B(n_1272),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1269),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1334),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1269),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1369),
.B(n_1407),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1356),
.A2(n_1322),
.B(n_1325),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1366),
.Y(n_1427)
);

AO32x2_ASAP7_75t_L g1428 ( 
.A1(n_1350),
.A2(n_1398),
.A3(n_1383),
.B1(n_1423),
.B2(n_1404),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1400),
.B(n_1235),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1356),
.A2(n_1261),
.B(n_1225),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1380),
.B(n_1238),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1378),
.A2(n_1231),
.B1(n_1339),
.B2(n_1329),
.C(n_1225),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1403),
.A2(n_1339),
.B(n_1329),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1405),
.A2(n_1332),
.B(n_1238),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_1236),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1405),
.A2(n_1236),
.B(n_1320),
.C(n_1223),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1359),
.A2(n_1223),
.B(n_1320),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1345),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1385),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1354),
.Y(n_1440)
);

OAI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1416),
.A2(n_1310),
.B(n_1317),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1389),
.B(n_1230),
.Y(n_1442)
);

OAI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1317),
.B(n_1335),
.C(n_1336),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1380),
.B(n_1390),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1389),
.B(n_1315),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1402),
.A2(n_1410),
.B(n_1413),
.C(n_1381),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1353),
.B(n_1390),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1410),
.A2(n_1344),
.B(n_1408),
.C(n_1401),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1393),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1410),
.A2(n_1344),
.B1(n_1408),
.B2(n_1401),
.C(n_1392),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_SL g1451 ( 
.A(n_1374),
.B(n_1420),
.Y(n_1451)
);

AOI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1392),
.A2(n_1394),
.B1(n_1365),
.B2(n_1367),
.C(n_1388),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1391),
.B(n_1384),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1398),
.B(n_1397),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1365),
.B(n_1367),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1403),
.A2(n_1411),
.B(n_1359),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1373),
.A2(n_1363),
.B(n_1349),
.C(n_1348),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1403),
.A2(n_1411),
.B(n_1399),
.Y(n_1458)
);

OAI21xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1422),
.A2(n_1424),
.B(n_1423),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1364),
.B(n_1418),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1355),
.B(n_1352),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1372),
.A2(n_1411),
.B(n_1370),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1411),
.A2(n_1387),
.B(n_1414),
.C(n_1386),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1412),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1399),
.A2(n_1409),
.B(n_1419),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1406),
.B(n_1395),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1415),
.Y(n_1467)
);

NOR3xp33_ASAP7_75t_SL g1468 ( 
.A(n_1421),
.B(n_1417),
.C(n_1419),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1406),
.B(n_1395),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1355),
.B(n_1352),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1362),
.Y(n_1471)
);

AO32x2_ASAP7_75t_L g1472 ( 
.A1(n_1404),
.A2(n_1362),
.A3(n_1396),
.B1(n_1368),
.B2(n_1371),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1427),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1472),
.B(n_1372),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1472),
.B(n_1372),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1472),
.B(n_1372),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1471),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.B(n_1362),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1425),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1426),
.A2(n_1414),
.B1(n_1379),
.B2(n_1357),
.Y(n_1480)
);

OR2x6_ASAP7_75t_SL g1481 ( 
.A(n_1435),
.B(n_1376),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1362),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1466),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1426),
.A2(n_1414),
.B1(n_1357),
.B2(n_1361),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_1461),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1438),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1428),
.B(n_1447),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1428),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1428),
.B(n_1375),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1461),
.B(n_1358),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1360),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1450),
.A2(n_1346),
.B1(n_1347),
.B2(n_1351),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1470),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1382),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1459),
.B(n_1395),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1494),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1490),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1480),
.A2(n_1446),
.B1(n_1463),
.B2(n_1448),
.C(n_1458),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1494),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1477),
.Y(n_1500)
);

OAI321xp33_ASAP7_75t_L g1501 ( 
.A1(n_1480),
.A2(n_1463),
.A3(n_1458),
.B1(n_1462),
.B2(n_1465),
.C(n_1434),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1474),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1490),
.Y(n_1503)
);

OAI33xp33_ASAP7_75t_L g1504 ( 
.A1(n_1478),
.A2(n_1435),
.A3(n_1441),
.B1(n_1445),
.B2(n_1442),
.B3(n_1429),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1487),
.B(n_1453),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1491),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1453),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1487),
.B(n_1467),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1487),
.B(n_1469),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1491),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1444),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1482),
.B(n_1437),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1464),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1492),
.A2(n_1452),
.B1(n_1434),
.B2(n_1432),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1454),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1473),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1486),
.B(n_1451),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1473),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1484),
.A2(n_1377),
.B1(n_1376),
.B2(n_1465),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1492),
.A2(n_1432),
.B1(n_1430),
.B2(n_1433),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1488),
.B(n_1444),
.Y(n_1523)
);

OAI31xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1495),
.A2(n_1430),
.A3(n_1443),
.B(n_1431),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1485),
.B(n_1457),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1518),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1517),
.B(n_1488),
.Y(n_1528)
);

AND2x4_ASAP7_75t_SL g1529 ( 
.A(n_1512),
.B(n_1468),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1517),
.B(n_1489),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1497),
.B(n_1493),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1518),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

AND2x2_ASAP7_75t_SL g1534 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1520),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1517),
.B(n_1489),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1526),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1506),
.Y(n_1538)
);

NAND2x1_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1525),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1513),
.B(n_1481),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1481),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1509),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1526),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1514),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1483),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1523),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1534),
.B(n_1524),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1523),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1544),
.B(n_1512),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1534),
.A2(n_1515),
.B1(n_1522),
.B2(n_1498),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1534),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1539),
.A2(n_1515),
.B1(n_1522),
.B2(n_1498),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1545),
.B(n_1508),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1549),
.B(n_1440),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1529),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1533),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1529),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1545),
.B(n_1508),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1499),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1535),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1529),
.B(n_1504),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1547),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1499),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1540),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1541),
.B(n_1542),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1541),
.A2(n_1443),
.B(n_1436),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1550),
.B(n_1500),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1554),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1552),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1576),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1581),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1581),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1576),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_L g1598 ( 
.A(n_1574),
.B(n_1542),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1562),
.B(n_1591),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1588),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1591),
.B(n_1554),
.Y(n_1602)
);

AOI211xp5_ASAP7_75t_L g1603 ( 
.A1(n_1564),
.A2(n_1570),
.B(n_1555),
.C(n_1582),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1563),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1560),
.B(n_1542),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1560),
.B(n_1543),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1543),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1564),
.B(n_1528),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1588),
.B(n_1543),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1563),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1557),
.B(n_1528),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1528),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1567),
.B(n_1521),
.C(n_1476),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1574),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1557),
.B(n_1553),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1566),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1566),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1551),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_L g1620 ( 
.A(n_1574),
.B(n_1460),
.C(n_1536),
.D(n_1530),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1567),
.A2(n_1501),
.B(n_1475),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1565),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1565),
.B(n_1551),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1568),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1603),
.A2(n_1567),
.B(n_1501),
.Y(n_1627)
);

OAI21xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1613),
.A2(n_1559),
.B(n_1536),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1604),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1584),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1604),
.Y(n_1631)
);

AOI211xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1598),
.A2(n_1584),
.B(n_1559),
.C(n_1578),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1622),
.A2(n_1589),
.B1(n_1539),
.B2(n_1476),
.C(n_1474),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1617),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1584),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1618),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1609),
.B(n_1559),
.Y(n_1638)
);

AOI222xp33_ASAP7_75t_L g1639 ( 
.A1(n_1614),
.A2(n_1475),
.B1(n_1476),
.B2(n_1504),
.C1(n_1502),
.C2(n_1530),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1589),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1623),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1626),
.Y(n_1642)
);

INVxp33_ASAP7_75t_L g1643 ( 
.A(n_1623),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1623),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1612),
.A2(n_1475),
.B(n_1476),
.C(n_1599),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1602),
.A2(n_1578),
.B(n_1580),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1600),
.B(n_1551),
.Y(n_1647)
);

NAND4xp25_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1571),
.C(n_1572),
.D(n_1577),
.Y(n_1648)
);

OAI21xp33_ASAP7_75t_L g1649 ( 
.A1(n_1620),
.A2(n_1572),
.B(n_1565),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1616),
.A2(n_1475),
.B1(n_1502),
.B2(n_1530),
.C(n_1536),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1615),
.A2(n_1580),
.B(n_1590),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1648),
.B(n_1638),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1629),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1630),
.B(n_1600),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1641),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1631),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1636),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1635),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1643),
.B(n_1610),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1640),
.B(n_1615),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1627),
.A2(n_1619),
.B(n_1605),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1643),
.Y(n_1665)
);

AOI222xp33_ASAP7_75t_L g1666 ( 
.A1(n_1645),
.A2(n_1633),
.B1(n_1628),
.B2(n_1650),
.C1(n_1637),
.C2(n_1642),
.Y(n_1666)
);

O2A1O1Ixp33_ASAP7_75t_SL g1667 ( 
.A1(n_1651),
.A2(n_1596),
.B(n_1595),
.C(n_1601),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1619),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1645),
.A2(n_1601),
.B(n_1593),
.Y(n_1669)
);

OAI322xp33_ASAP7_75t_L g1670 ( 
.A1(n_1647),
.A2(n_1593),
.A3(n_1612),
.B1(n_1592),
.B2(n_1624),
.C1(n_1621),
.C2(n_1569),
.Y(n_1670)
);

AO22x2_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1661),
.B1(n_1653),
.B2(n_1656),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1662),
.B(n_1606),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1665),
.B(n_1660),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1658),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1657),
.B(n_1608),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1649),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1663),
.Y(n_1678)
);

XNOR2x1_ASAP7_75t_L g1679 ( 
.A(n_1658),
.B(n_1652),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1655),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1655),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1673),
.B(n_1668),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1673),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1674),
.A2(n_1669),
.B(n_1664),
.C(n_1665),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1676),
.B(n_1657),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1678),
.A2(n_1667),
.B(n_1670),
.C(n_1666),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_1667),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1671),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1671),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1671),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_SL g1691 ( 
.A(n_1672),
.B(n_1677),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1686),
.A2(n_1675),
.B1(n_1681),
.B2(n_1680),
.C(n_1654),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1679),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1687),
.A2(n_1605),
.B(n_1639),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1685),
.B(n_1606),
.Y(n_1696)
);

AOI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1687),
.A2(n_1624),
.B(n_1621),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_L g1698 ( 
.A(n_1696),
.B(n_1683),
.Y(n_1698)
);

OAI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1694),
.A2(n_1690),
.B(n_1689),
.C(n_1682),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1692),
.A2(n_1691),
.B(n_1592),
.C(n_1575),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1693),
.A2(n_1478),
.B1(n_1575),
.B2(n_1556),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1697),
.A2(n_1625),
.B(n_1607),
.C(n_1579),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1695),
.A2(n_1579),
.B1(n_1585),
.B2(n_1556),
.C(n_1575),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1703),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1702),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1698),
.A2(n_1585),
.B1(n_1556),
.B2(n_1579),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1699),
.B(n_1607),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1700),
.Y(n_1708)
);

NAND3x1_ASAP7_75t_L g1709 ( 
.A(n_1708),
.B(n_1625),
.C(n_1571),
.Y(n_1709)
);

XOR2x2_ASAP7_75t_L g1710 ( 
.A(n_1707),
.B(n_1701),
.Y(n_1710)
);

OAI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1705),
.A2(n_1583),
.B(n_1585),
.C(n_1586),
.Y(n_1711)
);

XNOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1710),
.B(n_1706),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1712),
.Y(n_1713)
);

AND2x2_ASAP7_75t_SL g1714 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1713),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1715),
.B(n_1704),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1714),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1717),
.Y(n_1718)
);

AO21x2_ASAP7_75t_L g1719 ( 
.A1(n_1716),
.A2(n_1711),
.B(n_1709),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1583),
.B(n_1586),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1718),
.B(n_1719),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1721),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1718),
.B1(n_1583),
.B2(n_1586),
.C(n_1568),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1590),
.B(n_1587),
.Y(n_1724)
);


endmodule