module fake_jpeg_28755_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_20),
.B1(n_16),
.B2(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_34),
.B1(n_26),
.B2(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_16),
.B1(n_17),
.B2(n_14),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_33),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_34),
.B1(n_27),
.B2(n_30),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_24),
.A3(n_29),
.B1(n_36),
.B2(n_11),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_21),
.B1(n_36),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_58),
.B1(n_35),
.B2(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_47),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_44),
.B1(n_46),
.B2(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_50),
.B(n_56),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_66),
.C(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_0),
.C(n_1),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

OA21x2_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_50),
.B(n_14),
.Y(n_75)
);

OA21x2_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_42),
.B(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_82),
.Y(n_90)
);

OAI322xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_50),
.A3(n_65),
.B1(n_64),
.B2(n_60),
.C1(n_63),
.C2(n_5),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_85),
.C(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_35),
.B1(n_49),
.B2(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_40),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_1),
.B(n_2),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_2),
.B(n_3),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_3),
.B(n_4),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_77),
.C(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_78),
.C(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_72),
.B1(n_78),
.B2(n_82),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_81),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.C(n_95),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_3),
.B(n_5),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_104),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_7),
.Y(n_107)
);


endmodule