module fake_jpeg_6629_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx12_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_40),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_59),
.B1(n_63),
.B2(n_15),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_25),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_18),
.B1(n_15),
.B2(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_18),
.B1(n_29),
.B2(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_30),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_37),
.C(n_40),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_73),
.C(n_78),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_63),
.B1(n_51),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_60),
.B1(n_41),
.B2(n_36),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_40),
.C(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_33),
.C(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_36),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_R g113 ( 
.A(n_87),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_91),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_51),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_92),
.B1(n_102),
.B2(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_43),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_98),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_56),
.C(n_52),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_47),
.C(n_72),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_44),
.B(n_57),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_72),
.B(n_77),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_87),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_83),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_80),
.B1(n_60),
.B2(n_74),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_83),
.B(n_65),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_100),
.B1(n_94),
.B2(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_117),
.Y(n_132)
);

OA21x2_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_119),
.B(n_104),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_128),
.B(n_26),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_124),
.B1(n_122),
.B2(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_19),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_100),
.C(n_17),
.Y(n_134)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_93),
.B(n_85),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_135),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_143),
.C(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_95),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_42),
.B1(n_75),
.B2(n_29),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_116),
.B1(n_110),
.B2(n_30),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_17),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_75),
.C(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_147),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_27),
.B(n_19),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_42),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_119),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_86),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_17),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_30),
.C(n_26),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_119),
.A3(n_112),
.B1(n_108),
.B2(n_125),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_126),
.B(n_31),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_165),
.B(n_168),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_159),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_27),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_28),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_135),
.B1(n_26),
.B2(n_21),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_137),
.C(n_143),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_164),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_131),
.B1(n_151),
.B2(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_145),
.B1(n_134),
.B2(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_189),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_144),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_152),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_17),
.B(n_24),
.C(n_16),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_163),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_23),
.C(n_20),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_157),
.B(n_155),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_202),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_154),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_203),
.B1(n_177),
.B2(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_176),
.B(n_171),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_160),
.B1(n_165),
.B2(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_161),
.C(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_187),
.C(n_190),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_153),
.B1(n_166),
.B2(n_161),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_190),
.B1(n_28),
.B2(n_23),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_175),
.B1(n_191),
.B2(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_212),
.B1(n_195),
.B2(n_192),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_214),
.B1(n_218),
.B2(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_201),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_211),
.A2(n_216),
.B(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_42),
.C(n_28),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_42),
.B1(n_0),
.B2(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_193),
.C(n_197),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_2),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_216),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_234),
.B(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_210),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_5),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_3),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_240),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_4),
.B(n_5),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_6),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_233),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_6),
.C2(n_13),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_246),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_14),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_239),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_245),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_11),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_12),
.Y(n_252)
);


endmodule