module fake_jpeg_13707_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_53),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_40),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_50),
.B1(n_41),
.B2(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_77),
.B1(n_23),
.B2(n_10),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_8),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_80),
.B(n_81),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_66),
.C(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_62),
.B1(n_43),
.B2(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_21),
.B(n_32),
.C(n_31),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_5),
.B(n_6),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_91),
.B1(n_92),
.B2(n_9),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_11),
.C(n_15),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_81),
.B1(n_69),
.B2(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_26),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_16),
.C(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_28),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_83),
.B1(n_91),
.B2(n_84),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.C(n_97),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_93),
.B(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

AOI321xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_87),
.A3(n_102),
.B1(n_33),
.B2(n_29),
.C(n_30),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_102),
.Y(n_108)
);


endmodule