module real_jpeg_18812_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_373),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_0),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

NAND2x1_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_66),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

NAND2x1_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_5),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_5),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_7),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_7),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_7),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_8),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_8),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_8),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_8),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_8),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_8),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_8),
.B(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_10),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g175 ( 
.A(n_12),
.Y(n_175)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_152),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_151),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_19),
.B(n_128),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_82),
.C(n_107),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_20),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_56),
.C(n_75),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_21),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_33),
.C(n_41),
.Y(n_21)
);

XOR2x1_ASAP7_75t_L g273 ( 
.A(n_22),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_23),
.A2(n_31),
.B1(n_207),
.B2(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B(n_28),
.Y(n_23)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_26),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_24),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_91),
.C(n_94),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_24),
.A2(n_77),
.B1(n_91),
.B2(n_92),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_24),
.A2(n_77),
.B1(n_176),
.B2(n_230),
.Y(n_348)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_25),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_35),
.B(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_29),
.C(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_26),
.A2(n_35),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_26),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_26),
.A2(n_164),
.B1(n_292),
.B2(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_28),
.B(n_29),
.C(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_28),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_29),
.A2(n_32),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_29),
.A2(n_32),
.B1(n_214),
.B2(n_215),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_31),
.A2(n_207),
.B(n_301),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_62),
.C(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_33),
.B(n_41),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_35),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_35),
.A2(n_59),
.B1(n_165),
.B2(n_169),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_35),
.B(n_59),
.C(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_35),
.A2(n_165),
.B1(n_302),
.B2(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_37),
.B(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_37),
.B(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_43),
.A2(n_44),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_43),
.A2(n_44),
.B1(n_91),
.B2(n_92),
.Y(n_342)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_44),
.B(n_47),
.C(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_44),
.B(n_79),
.C(n_112),
.Y(n_134)
);

O2A1O1Ixp5_ASAP7_75t_L g200 ( 
.A1(n_44),
.A2(n_92),
.B(n_201),
.C(n_206),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_45),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_52),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_52),
.A2(n_123),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_52),
.A2(n_65),
.B1(n_123),
.B2(n_145),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_52),
.B(n_145),
.C(n_289),
.Y(n_313)
);

OR2x4_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_54),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_95),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_55),
.B(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_56),
.B(n_75),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.C(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_57),
.A2(n_58),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.C(n_65),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_59),
.A2(n_65),
.B1(n_145),
.B2(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_59),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_86),
.B1(n_87),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_62),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_62),
.A2(n_127),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_62),
.B(n_72),
.C(n_240),
.Y(n_346)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_65),
.A2(n_101),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_65),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_65),
.A2(n_147),
.B(n_148),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_65),
.B(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_68),
.B(n_72),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_68),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_69),
.B(n_172),
.C(n_176),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_72),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

AOI22x1_ASAP7_75t_SL g244 ( 
.A1(n_71),
.A2(n_72),
.B1(n_179),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_76),
.C(n_79),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_72),
.B(n_171),
.C(n_179),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_72),
.B(n_196),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_74),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_77),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_81),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_79),
.B(n_92),
.C(n_101),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_79),
.A2(n_81),
.B1(n_100),
.B2(n_105),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_82),
.B(n_107),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_99),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_90),
.C(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_91),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_91),
.B(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_91),
.B(n_325),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_119),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_94),
.B(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_94),
.A2(n_232),
.B(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_101),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_103),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_101),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_101),
.A2(n_144),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_101),
.A2(n_206),
.B(n_207),
.C(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_101),
.A2(n_144),
.B1(n_207),
.B2(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_116),
.C(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_124),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_124),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_123),
.B(n_212),
.C(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_150),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_140),
.B1(n_141),
.B2(n_149),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_187),
.B(n_371),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_185),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_154),
.B(n_185),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_R g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_155),
.B(n_157),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_159),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_170),
.C(n_181),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_160),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.C(n_167),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_167),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_170),
.A2(n_181),
.B1(n_182),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_172),
.A2(n_176),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI321xp33_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_264),
.A3(n_281),
.B1(n_364),
.B2(n_365),
.C(n_370),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI31xp33_ASAP7_75t_L g365 ( 
.A1(n_190),
.A2(n_277),
.A3(n_366),
.B(n_369),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_253),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_191),
.B(n_253),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_223),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_192),
.B(n_224),
.C(n_249),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_211),
.C(n_219),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_199),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_194),
.B(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_198),
.B(n_200),
.Y(n_356)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_201),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_201),
.A2(n_289),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_219),
.B1(n_220),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_248),
.B2(n_249),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_241),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.C(n_239),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_230),
.B(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_230),
.A2(n_291),
.B(n_292),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_232),
.B1(n_239),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_271),
.C(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_254),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_257),
.B(n_260),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_261),
.B(n_263),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_262),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_277),
.Y(n_264)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_265),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_266),
.B(n_275),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.C(n_273),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_273),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_278),
.B(n_280),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_360),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_350),
.B(n_359),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_333),
.B(n_349),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_314),
.B(n_332),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_298),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_295),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_307),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_308),
.C(n_313),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_324),
.B(n_326),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_322),
.B(n_331),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_319),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_327),
.B(n_330),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_335),
.Y(n_349)
);

XOR2x2_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_339),
.C(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_345),
.C(n_348),
.Y(n_354)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_355),
.C(n_357),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_362),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);


endmodule