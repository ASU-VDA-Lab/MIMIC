module fake_jpeg_14132_n_91 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx11_ASAP7_75t_SL g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_8),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_0),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_10),
.B(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_21),
.C(n_20),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_41),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI22x1_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_55),
.B(n_46),
.C(n_49),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_54),
.B(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_29),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_12),
.B1(n_10),
.B2(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_54),
.C(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_61),
.B1(n_1),
.B2(n_4),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_37),
.B1(n_39),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_37),
.B1(n_23),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_52),
.B(n_53),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_52),
.B1(n_48),
.B2(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_69),
.B1(n_63),
.B2(n_64),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_68),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_71),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_46),
.B(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.C(n_64),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.C(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_65),
.C(n_71),
.Y(n_79)
);

AOI21x1_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_83),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_5),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_6),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_74),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_69),
.B(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_6),
.Y(n_91)
);


endmodule