module fake_jpeg_20458_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_27),
.B1(n_15),
.B2(n_13),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_63),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_34),
.B1(n_48),
.B2(n_45),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_61),
.A2(n_78),
.B1(n_88),
.B2(n_16),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_19),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_67),
.C(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_66),
.B1(n_74),
.B2(n_79),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_65),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_36),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_71),
.B(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_22),
.B1(n_29),
.B2(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_75),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_18),
.B1(n_30),
.B2(n_31),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_57),
.B1(n_49),
.B2(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_14),
.B1(n_31),
.B2(n_38),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_30),
.B1(n_15),
.B2(n_13),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_90),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_14),
.B1(n_42),
.B2(n_21),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_92),
.B1(n_13),
.B2(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_93),
.Y(n_113)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_14),
.B1(n_23),
.B2(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_17),
.A3(n_20),
.B1(n_40),
.B2(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_11),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_51),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_117),
.B1(n_132),
.B2(n_85),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_112),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_16),
.C(n_26),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_60),
.B1(n_70),
.B2(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_16),
.B1(n_26),
.B2(n_2),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_158),
.B1(n_124),
.B2(n_126),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_80),
.B1(n_76),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_138),
.B1(n_150),
.B2(n_157),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_62),
.B1(n_64),
.B2(n_77),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_145),
.B(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_140),
.Y(n_173)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_126),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_107),
.C(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_151),
.C(n_104),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_101),
.B(n_119),
.C(n_120),
.D(n_123),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_109),
.C(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_16),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_148),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_16),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_89),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_87),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_72),
.B1(n_73),
.B2(n_94),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_86),
.C(n_12),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_11),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_104),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_141),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_116),
.C(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_135),
.C(n_142),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_131),
.Y(n_166)
);

OAI22x1_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_105),
.B1(n_132),
.B2(n_130),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_175),
.B1(n_179),
.B2(n_145),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_124),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_171),
.B(n_129),
.Y(n_203)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_1),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_109),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_183),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_115),
.B1(n_108),
.B2(n_129),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_187),
.C(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_197),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_147),
.B(n_139),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_168),
.B(n_166),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_140),
.B1(n_157),
.B2(n_158),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_193),
.B1(n_175),
.B2(n_179),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_153),
.B1(n_155),
.B2(n_122),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_145),
.C(n_122),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_205),
.B1(n_163),
.B2(n_178),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_109),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_201),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_110),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_110),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_207),
.B(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_5),
.C(n_6),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_210),
.A2(n_221),
.B(n_225),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_190),
.B1(n_203),
.B2(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_223),
.B1(n_199),
.B2(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_222),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_172),
.B(n_171),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_182),
.C(n_162),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_169),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_187),
.C(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_229),
.C(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_208),
.C(n_196),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_209),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_236),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_204),
.C(n_193),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_192),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_201),
.C(n_197),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_188),
.B(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_184),
.C(n_170),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_254),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_225),
.B1(n_215),
.B2(n_220),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_255),
.B(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_242),
.C(n_235),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_265),
.C(n_248),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_244),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_244),
.B(n_233),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_236),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_238),
.C(n_239),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_271),
.B(n_272),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_260),
.A2(n_259),
.B(n_258),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_270),
.A3(n_261),
.B1(n_263),
.B2(n_200),
.C1(n_264),
.C2(n_184),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_247),
.C(n_217),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_274),
.B(n_8),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_200),
.A3(n_170),
.B1(n_261),
.B2(n_220),
.C1(n_180),
.C2(n_6),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_7),
.C(n_8),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_271),
.B1(n_267),
.B2(n_9),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_279),
.C(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_9),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_9),
.C(n_10),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_10),
.Y(n_284)
);


endmodule