module fake_jpeg_4541_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_39),
.B1(n_19),
.B2(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_25),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_21),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_54),
.B1(n_59),
.B2(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_25),
.C(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_26),
.B1(n_33),
.B2(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_29),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_72),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_85),
.B1(n_66),
.B2(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_56),
.A3(n_55),
.B1(n_68),
.B2(n_67),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_90),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_43),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_94),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_68),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_101),
.B1(n_82),
.B2(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_53),
.B(n_60),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_28),
.A3(n_43),
.B1(n_17),
.B2(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_51),
.B1(n_54),
.B2(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_32),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_38),
.B1(n_21),
.B2(n_17),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_40),
.C(n_65),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_97),
.C(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_39),
.B1(n_40),
.B2(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_69),
.B(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_124),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_66),
.B1(n_43),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_76),
.B1(n_95),
.B2(n_71),
.Y(n_160)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_90),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_92),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_42),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_115),
.C(n_114),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_134),
.A2(n_157),
.B(n_24),
.Y(n_186)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_140),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_88),
.B1(n_105),
.B2(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_160),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_81),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_81),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_89),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_89),
.B1(n_87),
.B2(n_99),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_152),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_103),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_102),
.B(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_107),
.Y(n_157)
);

OAI22x1_ASAP7_75t_L g158 ( 
.A1(n_110),
.A2(n_73),
.B1(n_87),
.B2(n_43),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_106),
.B1(n_121),
.B2(n_116),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_72),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_102),
.A2(n_73),
.B1(n_70),
.B2(n_79),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_34),
.B1(n_24),
.B2(n_22),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_170),
.B(n_182),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_164),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_180),
.C(n_188),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_120),
.B(n_128),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_167),
.B(n_177),
.CI(n_186),
.CON(n_203),
.SN(n_203)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_120),
.B(n_116),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_174),
.B1(n_178),
.B2(n_194),
.Y(n_218)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_121),
.B1(n_86),
.B2(n_43),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_42),
.B(n_29),
.C(n_24),
.D(n_22),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_34),
.B1(n_32),
.B2(n_42),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_163),
.B1(n_195),
.B2(n_171),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_42),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_193),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_24),
.A3(n_29),
.B1(n_78),
.B2(n_3),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_185),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_190),
.B1(n_149),
.B2(n_140),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_29),
.C(n_1),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_29),
.B(n_1),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_187),
.C(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_146),
.B1(n_139),
.B2(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_206),
.B1(n_215),
.B2(n_182),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_144),
.B1(n_133),
.B2(n_134),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_210),
.B(n_189),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_131),
.B(n_141),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_211),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_220),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_131),
.B1(n_161),
.B2(n_137),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_191),
.C(n_166),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_222),
.C(n_168),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_132),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_132),
.C(n_4),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_0),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_4),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_226),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_235),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_165),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_184),
.B1(n_167),
.B2(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_213),
.B1(n_218),
.B2(n_224),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_177),
.B1(n_164),
.B2(n_188),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_217),
.B(n_197),
.C(n_203),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_194),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_197),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_179),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_200),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_199),
.C(n_222),
.Y(n_272)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_218),
.B1(n_207),
.B2(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_8),
.B(n_9),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_249),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_260),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_223),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_264),
.B1(n_250),
.B2(n_247),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_271),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_242),
.B1(n_233),
.B2(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_267),
.C(n_272),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_270),
.B(n_229),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_232),
.B(n_203),
.Y(n_269)
);

BUFx12f_ASAP7_75t_SL g281 ( 
.A(n_269),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_199),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_202),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_235),
.C(n_228),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_277),
.C(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_238),
.C(n_239),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_234),
.B(n_231),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_265),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_251),
.B1(n_230),
.B2(n_246),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_288),
.B1(n_261),
.B2(n_198),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_286),
.B(n_264),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_261),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_240),
.B(n_243),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_230),
.B1(n_241),
.B2(n_237),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_241),
.C(n_198),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_262),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_262),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_304),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_267),
.C(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_301),
.C(n_288),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_269),
.B1(n_270),
.B2(n_252),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_280),
.B1(n_274),
.B2(n_11),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_275),
.B1(n_278),
.B2(n_284),
.C(n_282),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_279),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_261),
.C(n_203),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_10),
.Y(n_304)
);

NAND2x1_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_312),
.B(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_313),
.C(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_9),
.C(n_10),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_10),
.B(n_11),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_9),
.C(n_11),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_302),
.B(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_301),
.B(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_321),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_323),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_304),
.B(n_12),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_12),
.C(n_13),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_13),
.C(n_14),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_14),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.C(n_308),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_306),
.B(n_310),
.Y(n_329)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_316),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_308),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.A3(n_333),
.B1(n_327),
.B2(n_334),
.C1(n_317),
.C2(n_312),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_9),
.B(n_15),
.Y(n_339)
);


endmodule