module fake_jpeg_11926_n_595 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_595);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx11_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx3_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_61),
.Y(n_178)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_66),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_33),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_71),
.B(n_77),
.Y(n_147)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx6p67_ASAP7_75t_R g149 ( 
.A(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_33),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_88),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_94),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_34),
.B(n_15),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_113),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_100),
.B(n_111),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_43),
.B(n_1),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_119),
.Y(n_163)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

BUFx16f_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_117),
.Y(n_146)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_118),
.B(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_28),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_121),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_28),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_58),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_47),
.B1(n_42),
.B2(n_50),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_129),
.A2(n_133),
.B(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_63),
.C(n_85),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_187),
.C(n_39),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_64),
.A2(n_47),
.B1(n_44),
.B2(n_23),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_45),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_74),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_136),
.B(n_142),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_137),
.B(n_143),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_32),
.B1(n_50),
.B2(n_26),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_139),
.A2(n_36),
.B1(n_19),
.B2(n_30),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_44),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_74),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_151),
.B(n_152),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_172),
.B(n_189),
.Y(n_245)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

INVx11_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_76),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_183),
.B(n_3),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_69),
.B(n_58),
.C(n_51),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_23),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_116),
.B(n_44),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_202),
.Y(n_255)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_192),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_118),
.B(n_51),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_110),
.B(n_21),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_200),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_104),
.B(n_21),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_108),
.B(n_26),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_95),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_44),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_205),
.B(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_206),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_129),
.A2(n_124),
.B1(n_103),
.B2(n_102),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_207),
.A2(n_248),
.B1(n_148),
.B2(n_168),
.Y(n_312)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g284 ( 
.A(n_209),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_210),
.A2(n_231),
.B1(n_265),
.B2(n_166),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_218),
.Y(n_293)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_212),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_39),
.C(n_49),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_213),
.B(n_187),
.C(n_178),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_146),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_216),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_157),
.B(n_82),
.Y(n_218)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_220),
.Y(n_287)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_224),
.Y(n_329)
);

CKINVDCx9p33_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_228),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_67),
.B1(n_60),
.B2(n_81),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_49),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_240),
.Y(n_322)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_235),
.Y(n_314)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_184),
.A2(n_45),
.B1(n_36),
.B2(n_30),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_238),
.A2(n_268),
.B1(n_271),
.B2(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_127),
.B(n_101),
.Y(n_240)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_243),
.Y(n_330)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_133),
.A2(n_83),
.B1(n_28),
.B2(n_5),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_145),
.Y(n_253)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

INVx4_ASAP7_75t_SL g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_254),
.Y(n_323)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_149),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_257),
.Y(n_279)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_145),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_147),
.B(n_2),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_260),
.Y(n_289)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_144),
.B(n_3),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_154),
.B(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_262),
.B(n_264),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_160),
.B(n_5),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_263),
.B(n_270),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_158),
.B(n_5),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_195),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_164),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_267),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_272),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_149),
.B(n_5),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_184),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_167),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_198),
.A2(n_7),
.B(n_9),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_274),
.B(n_218),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_315),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_205),
.A2(n_125),
.B1(n_169),
.B2(n_132),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_286),
.A2(n_312),
.B1(n_162),
.B2(n_209),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_149),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_238),
.A2(n_181),
.B1(n_148),
.B2(n_131),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_297),
.B1(n_298),
.B2(n_305),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_217),
.A2(n_204),
.B1(n_177),
.B2(n_191),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_219),
.A2(n_186),
.B1(n_166),
.B2(n_181),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_248),
.A2(n_167),
.B1(n_159),
.B2(n_178),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_301),
.A2(n_325),
.B(n_194),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_156),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_249),
.C(n_230),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_231),
.A2(n_180),
.B1(n_203),
.B2(n_132),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_255),
.A2(n_203),
.B1(n_138),
.B2(n_155),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_320),
.A2(n_326),
.B1(n_224),
.B2(n_221),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_174),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_327),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_273),
.A2(n_168),
.B1(n_196),
.B2(n_194),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_138),
.B1(n_155),
.B2(n_162),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_251),
.B(n_180),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_233),
.B(n_229),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_322),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_297),
.A2(n_223),
.B(n_156),
.C(n_250),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_359),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_350),
.C(n_321),
.Y(n_392)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_289),
.B(n_216),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_340),
.B(n_343),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_223),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_347),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_214),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_345),
.B(n_279),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_236),
.Y(n_347)
);

INVx13_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_348),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_252),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_361),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_254),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_226),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_L g404 ( 
.A1(n_351),
.A2(n_354),
.B(n_355),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_324),
.B(n_325),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_281),
.B(n_309),
.Y(n_391)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_323),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_237),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_367),
.Y(n_394)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_301),
.A2(n_259),
.B1(n_250),
.B2(n_227),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_358),
.A2(n_362),
.B1(n_305),
.B2(n_291),
.Y(n_379)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_316),
.B(n_230),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_373),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_333),
.B(n_196),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_242),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_366),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_364),
.A2(n_285),
.B1(n_284),
.B2(n_310),
.Y(n_390)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_256),
.C(n_235),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_257),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_253),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_370),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_269),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_374),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_312),
.A2(n_228),
.B(n_267),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_299),
.Y(n_371)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_280),
.B(n_327),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_377),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_307),
.B(n_165),
.Y(n_374)
);

AOI22x1_ASAP7_75t_SL g375 ( 
.A1(n_298),
.A2(n_165),
.B1(n_246),
.B2(n_268),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_376),
.B(n_318),
.Y(n_412)
);

FAx1_ASAP7_75t_L g376 ( 
.A(n_288),
.B(n_164),
.CI(n_271),
.CON(n_376),
.SN(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_291),
.B(n_164),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_335),
.Y(n_421)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_393),
.B1(n_409),
.B2(n_414),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_391),
.A2(n_399),
.B(n_402),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_407),
.C(n_345),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_341),
.A2(n_336),
.B1(n_339),
.B2(n_352),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_346),
.A2(n_314),
.B(n_328),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_306),
.B1(n_319),
.B2(n_334),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_411),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_346),
.A2(n_287),
.B(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_405),
.Y(n_417)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_357),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_341),
.A2(n_339),
.B1(n_375),
.B2(n_372),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_336),
.A2(n_306),
.B1(n_334),
.B2(n_319),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_412),
.A2(n_354),
.B(n_376),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_376),
.A2(n_284),
.B1(n_308),
.B2(n_330),
.Y(n_414)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_399),
.A2(n_412),
.B(n_402),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_420),
.A2(n_424),
.B(n_437),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_421),
.A2(n_444),
.B1(n_300),
.B2(n_296),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_422),
.B(n_436),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_423),
.A2(n_447),
.B(n_424),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_381),
.A2(n_373),
.B(n_354),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_360),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_359),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_392),
.B(n_350),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_427),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_435),
.C(n_403),
.Y(n_457)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_396),
.A3(n_413),
.B1(n_393),
.B2(n_394),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_438),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_396),
.B1(n_410),
.B2(n_385),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_445),
.B(n_388),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_356),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_431),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_368),
.Y(n_432)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_351),
.C(n_355),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_401),
.Y(n_436)
);

AOI21xp33_ASAP7_75t_SL g437 ( 
.A1(n_381),
.A2(n_351),
.B(n_342),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_382),
.B(n_367),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_335),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_420),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_380),
.B(n_330),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_440),
.B(n_441),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_371),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_446),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_383),
.B(n_370),
.Y(n_443)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_408),
.A2(n_364),
.B(n_370),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_413),
.A2(n_377),
.B(n_332),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_300),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_318),
.B(n_317),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_411),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_SL g476 ( 
.A(n_449),
.B(n_348),
.C(n_329),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_451),
.A2(n_453),
.B(n_462),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_400),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_379),
.B1(n_408),
.B2(n_389),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_470),
.B1(n_444),
.B2(n_421),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_463),
.C(n_477),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_459),
.A2(n_472),
.B1(n_443),
.B2(n_431),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_418),
.A2(n_387),
.B(n_406),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_387),
.C(n_385),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_418),
.A2(n_415),
.B(n_405),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_447),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_384),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_428),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_397),
.B1(n_415),
.B2(n_384),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_417),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_471),
.B(n_474),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_478),
.B1(n_416),
.B2(n_449),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_417),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_476),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_294),
.C(n_317),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_292),
.B1(n_296),
.B2(n_311),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_425),
.B(n_311),
.Y(n_479)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_479),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_437),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_483),
.B(n_501),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_432),
.C(n_439),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_469),
.C(n_477),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_486),
.Y(n_511)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_488),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_503),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_493),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_438),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_491),
.B(n_498),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_492),
.A2(n_478),
.B1(n_453),
.B2(n_467),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_464),
.B1(n_459),
.B2(n_466),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_496),
.Y(n_522)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_441),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_497),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_436),
.Y(n_498)
);

BUFx4f_ASAP7_75t_SL g499 ( 
.A(n_450),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_458),
.B(n_419),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_462),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_439),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_470),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_455),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_505),
.B(n_463),
.Y(n_507)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_507),
.Y(n_529)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_500),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_513),
.A2(n_524),
.B(n_451),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_468),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_517),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_516),
.B(n_519),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_481),
.B(n_466),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_482),
.B(n_450),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_520),
.B(n_525),
.Y(n_531)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_523),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_492),
.A2(n_451),
.B(n_421),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_433),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_468),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_515),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_510),
.A2(n_480),
.B1(n_504),
.B2(n_494),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_528),
.A2(n_541),
.B1(n_543),
.B2(n_524),
.Y(n_557)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_534),
.B(n_444),
.Y(n_559)
);

A2O1A1O1Ixp25_ASAP7_75t_L g535 ( 
.A1(n_513),
.A2(n_502),
.B(n_484),
.C(n_501),
.D(n_496),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_535),
.A2(n_521),
.B(n_517),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_506),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_482),
.C(n_503),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_538),
.B(n_539),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_502),
.C(n_483),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_493),
.Y(n_542)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_542),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_518),
.A2(n_526),
.B1(n_486),
.B2(n_480),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_497),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_545),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_490),
.C(n_416),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_547),
.B(n_549),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_509),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_553),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_506),
.Y(n_549)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_550),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_518),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_524),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_554),
.B(n_448),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_545),
.C(n_533),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_555),
.B(n_558),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_510),
.Y(n_556)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_557),
.B(n_559),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_508),
.C(n_429),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_555),
.B(n_537),
.C(n_530),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_562),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_539),
.C(n_534),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_556),
.B(n_512),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_563),
.A2(n_440),
.B(n_558),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_560),
.A2(n_529),
.B1(n_531),
.B2(n_543),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_569),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_559),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_564),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_572),
.B(n_575),
.Y(n_582)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_554),
.Y(n_573)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_573),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_551),
.C(n_552),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_576),
.B(n_577),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_508),
.B1(n_559),
.B2(n_448),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_578),
.A2(n_565),
.B1(n_429),
.B2(n_549),
.Y(n_581)
);

AOI221xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_565),
.B1(n_570),
.B2(n_562),
.C(n_547),
.Y(n_580)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_580),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_581),
.B(n_572),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_574),
.A2(n_568),
.B(n_499),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_584),
.A2(n_573),
.B(n_446),
.Y(n_588)
);

NOR4xp25_ASAP7_75t_L g589 ( 
.A(n_587),
.B(n_582),
.C(n_580),
.D(n_585),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_586),
.C(n_583),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_589),
.A2(n_590),
.B(n_499),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_591),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_592),
.A2(n_294),
.B(n_292),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_277),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_277),
.Y(n_595)
);


endmodule