module fake_jpeg_6818_n_233 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_21),
.B1(n_16),
.B2(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_21),
.B1(n_25),
.B2(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_33),
.B1(n_25),
.B2(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_48),
.B1(n_39),
.B2(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_68),
.Y(n_85)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_13),
.B1(n_26),
.B2(n_23),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_29),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_71),
.B1(n_73),
.B2(n_59),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_40),
.B1(n_45),
.B2(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_40),
.B1(n_31),
.B2(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx24_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_66),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_52),
.B(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_56),
.B1(n_40),
.B2(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_85),
.B1(n_73),
.B2(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_95),
.B1(n_103),
.B2(n_105),
.Y(n_121)
);

INVxp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_68),
.C(n_31),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_50),
.C(n_35),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_10),
.Y(n_100)
);

XOR2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_57),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_22),
.B(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_50),
.B1(n_42),
.B2(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_72),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_27),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_84),
.B1(n_85),
.B2(n_69),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_117),
.B1(n_122),
.B2(n_124),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_86),
.B1(n_88),
.B2(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_118),
.B1(n_126),
.B2(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_120),
.B1(n_125),
.B2(n_119),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_35),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_123),
.C(n_30),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_56),
.B1(n_88),
.B2(n_65),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_56),
.B1(n_63),
.B2(n_51),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_30),
.B(n_27),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_51),
.B1(n_70),
.B2(n_72),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_79),
.B1(n_30),
.B2(n_27),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_64),
.B1(n_53),
.B2(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_102),
.A3(n_103),
.B1(n_94),
.B2(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_137),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_136),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_100),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_133),
.B(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.C(n_118),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_35),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_96),
.B1(n_79),
.B2(n_53),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_114),
.B1(n_81),
.B2(n_14),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_96),
.B1(n_81),
.B2(n_14),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_64),
.B1(n_19),
.B2(n_18),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_128),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_156),
.C(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_115),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_110),
.C(n_109),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_109),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_145),
.B1(n_132),
.B2(n_19),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_164),
.B1(n_132),
.B2(n_19),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_57),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_135),
.B(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_172),
.C(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_171),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_133),
.C(n_134),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_161),
.Y(n_174)
);

AO221x1_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_151),
.B1(n_165),
.B2(n_159),
.C(n_163),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_158),
.CI(n_162),
.CON(n_186),
.SN(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_57),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_20),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_154),
.C(n_160),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_18),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_158),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_193),
.C(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_192),
.B(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_150),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_197),
.C(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_190),
.B1(n_184),
.B2(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_152),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_202),
.B(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_168),
.C(n_8),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_8),
.C(n_12),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_205),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_188),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_186),
.B1(n_185),
.B2(n_184),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_5),
.B(n_10),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_18),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_4),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_14),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_205),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_214),
.B(n_215),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_4),
.B(n_9),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_212),
.A2(n_4),
.B(n_7),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_5),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_209),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_224),
.B(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_207),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_226),
.B(n_227),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_223),
.C(n_11),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_228),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_232),
.B(n_0),
.CI(n_1),
.CON(n_233),
.SN(n_233)
);


endmodule