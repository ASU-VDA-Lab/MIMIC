module fake_jpeg_16886_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_33),
.B(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_12),
.B(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_36),
.B1(n_18),
.B2(n_17),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_41),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_42),
.B(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_52),
.B(n_23),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_32),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_13),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_43),
.B1(n_29),
.B2(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_40),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_74),
.B1(n_67),
.B2(n_57),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_43),
.B1(n_29),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_69),
.B1(n_74),
.B2(n_72),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_59),
.C(n_49),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.C(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_51),
.C(n_46),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_84),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_54),
.C(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_63),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_67),
.B(n_61),
.C(n_48),
.D(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_98),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_91),
.C(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_76),
.B(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_102),
.B(n_25),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_77),
.C(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_64),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_99),
.A3(n_95),
.B1(n_96),
.B2(n_71),
.C1(n_13),
.C2(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_108),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_8),
.B(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_10),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_8),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_1),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_2),
.C(n_3),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C(n_111),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_13),
.C(n_5),
.Y(n_115)
);


endmodule