module fake_jpeg_8414_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_42),
.C(n_22),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.C(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_60),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_16),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_30),
.B1(n_29),
.B2(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_37),
.B1(n_34),
.B2(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_37),
.B1(n_34),
.B2(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_69),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_35),
.B(n_42),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_36),
.B1(n_41),
.B2(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_29),
.B1(n_17),
.B2(n_19),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_80),
.B(n_20),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_19),
.B1(n_17),
.B2(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

AOI22x1_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_35),
.B1(n_42),
.B2(n_36),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_35),
.B1(n_33),
.B2(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_36),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_96),
.B(n_111),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_40),
.C(n_39),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.C(n_103),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_69),
.B1(n_67),
.B2(n_75),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_41),
.B1(n_55),
.B2(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_104),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_64),
.C(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_27),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_41),
.B1(n_40),
.B2(n_16),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_56),
.B1(n_39),
.B2(n_40),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_40),
.B1(n_39),
.B2(n_18),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_63),
.B1(n_81),
.B2(n_76),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_86),
.B(n_39),
.C(n_26),
.D(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_135),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_124),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_134),
.B1(n_113),
.B2(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_106),
.C(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_78),
.B1(n_61),
.B2(n_47),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_78),
.B1(n_107),
.B2(n_43),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_61),
.C(n_1),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_32),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_100),
.B1(n_97),
.B2(n_89),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_150),
.B1(n_152),
.B2(n_158),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_89),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_98),
.B1(n_92),
.B2(n_95),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_24),
.B(n_4),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_118),
.B1(n_32),
.B2(n_24),
.C(n_5),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_43),
.C(n_83),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_78),
.B1(n_107),
.B2(n_47),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_161),
.B(n_162),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_116),
.B1(n_131),
.B2(n_119),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_0),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_144),
.B(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_26),
.B1(n_32),
.B2(n_25),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_32),
.B1(n_25),
.B2(n_83),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_114),
.B1(n_128),
.B2(n_112),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_32),
.B1(n_24),
.B2(n_0),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_177),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_182),
.B(n_162),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_24),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_24),
.C(n_6),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_2),
.C(n_6),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_2),
.C(n_9),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_149),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_9),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_155),
.C(n_160),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_138),
.C(n_139),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_9),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_187),
.B(n_193),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_144),
.B(n_142),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_191),
.B(n_182),
.Y(n_202)
);

OA21x2_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_156),
.B(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_142),
.B1(n_158),
.B2(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_184),
.B1(n_188),
.B2(n_171),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_151),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_165),
.C(n_176),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_206),
.C(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_170),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_164),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_212),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_164),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.C(n_169),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_153),
.Y(n_212)
);

OAI21x1_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_186),
.B(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_190),
.B(n_192),
.C(n_171),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_159),
.B(n_11),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_195),
.B1(n_191),
.B2(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_159),
.B1(n_197),
.B2(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_216),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_218),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_10),
.C(n_11),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_210),
.B1(n_201),
.B2(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_228),
.B(n_231),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_223),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_231),
.C(n_227),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_229),
.C(n_224),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_236),
.B1(n_241),
.B2(n_12),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.C(n_13),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_13),
.B(n_242),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_13),
.Y(n_248)
);


endmodule