module fake_jpeg_2373_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_48),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_1),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_64),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_72),
.Y(n_137)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_3),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_4),
.C(n_5),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_80),
.B(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_32),
.B(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_11),
.Y(n_121)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_16),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_19),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_17),
.B1(n_37),
.B2(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_107),
.B1(n_109),
.B2(n_112),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_4),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_99),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_29),
.B1(n_37),
.B2(n_35),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_103),
.B(n_115),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_38),
.B1(n_34),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_38),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_106),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_128),
.B1(n_95),
.B2(n_135),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_10),
.B1(n_11),
.B2(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_90),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_134),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_50),
.A2(n_51),
.B1(n_70),
.B2(n_67),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_45),
.B1(n_68),
.B2(n_88),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_92),
.B1(n_97),
.B2(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_65),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_52),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_91),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_143),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_144),
.A2(n_176),
.B1(n_177),
.B2(n_172),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_162),
.B1(n_113),
.B2(n_100),
.Y(n_182)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_146),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_111),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_150),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_132),
.C(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_158),
.C(n_172),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_99),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_161),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_104),
.C(n_136),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_107),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_115),
.B(n_101),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_171),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_152),
.B1(n_171),
.B2(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_155),
.Y(n_196)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_115),
.B1(n_100),
.B2(n_125),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_182),
.B1(n_187),
.B2(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_130),
.B1(n_133),
.B2(n_131),
.Y(n_187)
);

NOR2x1_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_148),
.B1(n_141),
.B2(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_186),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_155),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_201),
.C(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_145),
.A2(n_173),
.B1(n_170),
.B2(n_140),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_146),
.A2(n_167),
.B1(n_169),
.B2(n_138),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_215),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_177),
.B1(n_188),
.B2(n_196),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_195),
.B1(n_192),
.B2(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_220),
.B1(n_208),
.B2(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_180),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_181),
.A2(n_194),
.B(n_186),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_200),
.B(n_185),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_224),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_178),
.Y(n_221)
);

NAND2x1_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_225),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_192),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_227),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_202),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_229),
.B(n_219),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_206),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_223),
.B1(n_224),
.B2(n_209),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_221),
.B1(n_225),
.B2(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_213),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_236),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_216),
.B1(n_209),
.B2(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_253),
.B1(n_255),
.B2(n_258),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_211),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_231),
.B1(n_246),
.B2(n_235),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_237),
.C(n_242),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_242),
.C(n_245),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_233),
.Y(n_269)
);

AOI31xp67_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_251),
.A3(n_235),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_230),
.B1(n_252),
.B2(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_277),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_233),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_231),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_255),
.B1(n_252),
.B2(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_278),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_238),
.B(n_236),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_236),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_261),
.B(n_238),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_236),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_264),
.C(n_254),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_284),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_276),
.B(n_275),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_263),
.B(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_287),
.B1(n_279),
.B2(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_290),
.B1(n_286),
.B2(n_263),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_288),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_273),
.C(n_232),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_278),
.C(n_232),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.C(n_239),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_261),
.Y(n_297)
);


endmodule