module fake_jpeg_28390_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_22),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_26),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_39),
.C(n_45),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_77),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_83),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_50),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_28),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_97),
.Y(n_108)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_31),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_89),
.B1(n_99),
.B2(n_100),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_20),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_23),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_39),
.C(n_43),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_34),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_40),
.B1(n_38),
.B2(n_22),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_60),
.B1(n_47),
.B2(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_44),
.A3(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_99),
.A3(n_100),
.B1(n_23),
.B2(n_96),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_126),
.B1(n_127),
.B2(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_59),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_105),
.B1(n_80),
.B2(n_71),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_82),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_30),
.B1(n_53),
.B2(n_68),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_103),
.B1(n_85),
.B2(n_93),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_75),
.B(n_11),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_75),
.B(n_104),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_138),
.A2(n_140),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_92),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_144),
.B(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_88),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_88),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_99),
.C(n_100),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_159),
.C(n_132),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_150),
.B1(n_117),
.B2(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_70),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_129),
.B(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_30),
.B1(n_27),
.B2(n_95),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_157),
.B(n_165),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_78),
.B1(n_71),
.B2(n_70),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_155),
.B1(n_12),
.B2(n_2),
.Y(n_203)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_80),
.C(n_68),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_74),
.B1(n_86),
.B2(n_82),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_163),
.B1(n_125),
.B2(n_128),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_34),
.B1(n_32),
.B2(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_102),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_113),
.B(n_14),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_102),
.Y(n_169)
);

XOR2x2_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_109),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_173),
.A2(n_176),
.B(n_201),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_194),
.C(n_160),
.Y(n_205)
);

XOR2x2_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_121),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_119),
.B(n_127),
.C(n_117),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_178),
.A2(n_3),
.B(n_4),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_179),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_162),
.B1(n_139),
.B2(n_148),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_114),
.B1(n_115),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_115),
.B1(n_133),
.B2(n_125),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_119),
.B1(n_107),
.B2(n_122),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_189),
.B1(n_191),
.B2(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_122),
.B1(n_131),
.B2(n_34),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_131),
.B1(n_34),
.B2(n_102),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_131),
.B1(n_32),
.B2(n_16),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_32),
.C(n_16),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_1),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_155),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_1),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_226),
.C(n_183),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_173),
.B(n_199),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_230),
.B(n_231),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_197),
.B(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_141),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_213),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_214),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_12),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_225),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_1),
.C(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_204),
.B1(n_218),
.B2(n_220),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_191),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_176),
.A2(n_3),
.B(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_202),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_207),
.B1(n_206),
.B2(n_212),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.C(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_171),
.C(n_172),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_181),
.B1(n_180),
.B2(n_201),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_247),
.B1(n_207),
.B2(n_229),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_194),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_201),
.B1(n_177),
.B2(n_189),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_200),
.B1(n_196),
.B2(n_190),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_204),
.B1(n_227),
.B2(n_225),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_190),
.C(n_178),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_211),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_196),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_256),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_177),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_262),
.C(n_270),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_249),
.C(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_269),
.Y(n_288)
);

AO22x1_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_209),
.B1(n_230),
.B2(n_215),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_216),
.C(n_214),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_251),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_235),
.B(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_266),
.A2(n_233),
.B(n_239),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_224),
.B1(n_219),
.B2(n_222),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_247),
.B1(n_244),
.B2(n_237),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_268),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_210),
.C(n_213),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_206),
.C(n_170),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_276),
.C(n_212),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_236),
.C(n_254),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_292),
.B1(n_5),
.B2(n_7),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_256),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_290),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_5),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_267),
.B1(n_262),
.B2(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_257),
.B1(n_274),
.B2(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_264),
.C(n_273),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_304),
.C(n_305),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_273),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_283),
.B(n_287),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_264),
.B1(n_261),
.B2(n_7),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_280),
.B1(n_279),
.B2(n_281),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_261),
.B1(n_6),
.B2(n_7),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_303),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_8),
.C(n_9),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_314),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_282),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_288),
.B1(n_8),
.B2(n_10),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_300),
.B1(n_305),
.B2(n_8),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_301),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_303),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_310),
.C(n_307),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_304),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_296),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_315),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_313),
.B(n_316),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_328),
.B(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_319),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_330),
.B(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_319),
.C(n_299),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_313),
.B1(n_329),
.B2(n_312),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_298),
.B(n_10),
.Y(n_337)
);


endmodule