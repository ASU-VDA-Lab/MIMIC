module real_jpeg_25830_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_2),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_39),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_2),
.B(n_51),
.C(n_53),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_108),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_2),
.B(n_66),
.C(n_79),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_2),
.A2(n_68),
.B(n_217),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_5),
.A2(n_44),
.B1(n_66),
.B2(n_67),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_84),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_28),
.B1(n_57),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_187)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_48),
.B1(n_66),
.B2(n_67),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_14),
.A2(n_27),
.B1(n_40),
.B2(n_42),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_14),
.A2(n_27),
.B1(n_66),
.B2(n_67),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_15),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_118),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_97),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_61),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_25),
.B(n_45),
.C(n_61),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_26),
.Y(n_99)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_28),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_32),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_32),
.A2(n_136),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_34),
.B(n_40),
.Y(n_117)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_35),
.A2(n_37),
.A3(n_42),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_38),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_38),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_42),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_40),
.B(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_43),
.Y(n_133)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_55),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_47),
.A2(n_49),
.B1(n_59),
.B2(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_49),
.A2(n_55),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_51),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_51),
.B(n_224),
.Y(n_223)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_106),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_59),
.A2(n_107),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_75),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_62),
.B(n_75),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_90),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_69),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_67),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_67),
.B(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_70),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_72),
.B(n_87),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_68),
.A2(n_69),
.B1(n_113),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_68),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_68),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_69),
.Y(n_230)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_73),
.B(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_74),
.B(n_156),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_76),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_76),
.A2(n_205),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_93),
.B1(n_94),
.B2(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_77),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_77),
.A2(n_94),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_82),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_81),
.A2(n_152),
.B(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_81),
.B(n_156),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_85),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_94),
.B(n_153),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_97),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.C(n_109),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_98),
.B(n_104),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_109),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_114),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_111),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_138),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_137),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_172),
.B(n_259),
.C(n_264),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_166),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.C(n_159),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_144),
.A2(n_145),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_150),
.C(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_158),
.B(n_159),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_253),
.B(n_258),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_206),
.B(n_252),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_195),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_195),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.C(n_192),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_181),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B(n_186),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_229),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_202),
.C(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_246),
.B(n_251),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_225),
.B(n_245),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_219),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_234),
.B(n_244),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_232),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_239),
.B(n_243),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);


endmodule