module fake_jpeg_29138_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_50),
.Y(n_117)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_72),
.Y(n_127)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_56),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_58),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_75),
.Y(n_118)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_0),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_15),
.B(n_1),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_18),
.B(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_82),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_16),
.B(n_3),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_17),
.Y(n_115)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_21),
.B1(n_40),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_89),
.A2(n_94),
.B1(n_101),
.B2(n_104),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_23),
.B1(n_22),
.B2(n_39),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_21),
.B1(n_40),
.B2(n_38),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_43),
.B1(n_34),
.B2(n_28),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_43),
.B1(n_34),
.B2(n_22),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_31),
.B1(n_35),
.B2(n_24),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_35),
.B1(n_31),
.B2(n_41),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_44),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_38),
.B1(n_26),
.B2(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_62),
.A2(n_33),
.B1(n_26),
.B2(n_31),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_49),
.A2(n_35),
.B1(n_24),
.B2(n_25),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_77),
.B1(n_56),
.B2(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_76),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_58),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_35),
.B1(n_25),
.B2(n_7),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_80),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_35),
.B1(n_25),
.B2(n_7),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_74),
.A2(n_25),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_136),
.B(n_169),
.Y(n_206)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_137),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_162),
.B(n_131),
.C(n_100),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_139),
.A2(n_146),
.B1(n_167),
.B2(n_103),
.Y(n_208)
);

OR2x2_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_72),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_140),
.B(n_142),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_141),
.B(n_143),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_86),
.A2(n_60),
.B1(n_46),
.B2(n_66),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_89),
.A2(n_61),
.B1(n_81),
.B2(n_73),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_45),
.B(n_64),
.C(n_85),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_163),
.C(n_172),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_79),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_111),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_149),
.Y(n_197)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_68),
.B1(n_45),
.B2(n_65),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_173),
.Y(n_220)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_52),
.B(n_47),
.C(n_8),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_52),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_170),
.Y(n_199)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_105),
.A2(n_103),
.B1(n_98),
.B2(n_129),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_R g163 ( 
.A(n_127),
.B(n_4),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_87),
.Y(n_166)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_167)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_117),
.B(n_9),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_10),
.Y(n_170)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_114),
.Y(n_172)
);

OR2x2_ASAP7_75t_SL g173 ( 
.A(n_109),
.B(n_104),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_112),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_179),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_11),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_14),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_12),
.B(n_13),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_13),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_102),
.C(n_100),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_101),
.A2(n_14),
.B1(n_92),
.B2(n_129),
.Y(n_181)
);

AO22x2_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_113),
.B1(n_102),
.B2(n_121),
.Y(n_186)
);

AO21x2_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_142),
.B(n_147),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_171),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_215),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_191),
.A2(n_14),
.B1(n_174),
.B2(n_212),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_108),
.C(n_90),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_214),
.C(n_188),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_218),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_161),
.B1(n_181),
.B2(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_150),
.B1(n_93),
.B2(n_164),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_137),
.B1(n_159),
.B2(n_91),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_125),
.B1(n_121),
.B2(n_88),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_151),
.B1(n_166),
.B2(n_149),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_108),
.C(n_133),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_88),
.B1(n_93),
.B2(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_148),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_230),
.B1(n_245),
.B2(n_251),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_248),
.B(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_180),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_170),
.B1(n_177),
.B2(n_140),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_179),
.B(n_156),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_216),
.B(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_238),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_233),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_241),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_235),
.Y(n_272)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_166),
.B(n_139),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_258),
.B1(n_208),
.B2(n_197),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_152),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_155),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_250),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_201),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_186),
.A2(n_119),
.B1(n_149),
.B2(n_168),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_204),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_222),
.C(n_210),
.Y(n_265)
);

OR2x4_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_132),
.Y(n_248)
);

XOR2x2_ASAP7_75t_SL g249 ( 
.A(n_214),
.B(n_91),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_259),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_174),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_183),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_196),
.Y(n_290)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_198),
.B(n_132),
.CI(n_174),
.CON(n_257),
.SN(n_257)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_212),
.B1(n_211),
.B2(n_190),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_260),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_185),
.C(n_209),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_274),
.C(n_275),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_257),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_282),
.B1(n_226),
.B2(n_250),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_218),
.B1(n_191),
.B2(n_205),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_270),
.A2(n_271),
.B1(n_286),
.B2(n_248),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_191),
.B1(n_197),
.B2(n_213),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_229),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_195),
.C(n_192),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_191),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_288),
.C(n_291),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_239),
.A2(n_213),
.B1(n_194),
.B2(n_184),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_194),
.B1(n_184),
.B2(n_187),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_221),
.C(n_196),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_300),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_277),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_235),
.B1(n_246),
.B2(n_237),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_317),
.B1(n_290),
.B2(n_260),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_272),
.B(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_309),
.B1(n_311),
.B2(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_307),
.B1(n_312),
.B2(n_296),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_224),
.B1(n_227),
.B2(n_242),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_257),
.B(n_234),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_316),
.B(n_280),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_227),
.B1(n_224),
.B2(n_254),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_227),
.B1(n_253),
.B2(n_238),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_228),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_236),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_319),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_283),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_283),
.C(n_274),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_322),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_263),
.C(n_262),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_263),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_334),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_287),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_336),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_327),
.A2(n_261),
.B(n_314),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_328),
.A2(n_330),
.B1(n_309),
.B2(n_303),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_269),
.C(n_267),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_338),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_306),
.A2(n_282),
.B1(n_271),
.B2(n_261),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_288),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_286),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_234),
.C(n_272),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_326),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_302),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_349),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_311),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_334),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_294),
.B(n_307),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_348),
.A2(n_321),
.B(n_328),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_300),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_350),
.A2(n_352),
.B(n_356),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_354),
.B1(n_357),
.B2(n_359),
.Y(n_367)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_321),
.A2(n_227),
.B(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_270),
.B1(n_295),
.B2(n_299),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_322),
.C(n_319),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_373),
.C(n_355),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_364),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_323),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_370),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_320),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_348),
.A2(n_358),
.B(n_342),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_372),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_369),
.A2(n_298),
.B(n_347),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_336),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_338),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_335),
.Y(n_373)
);

AOI322xp5_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_353),
.A3(n_352),
.B1(n_356),
.B2(n_295),
.C1(n_344),
.C2(n_349),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_377),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_367),
.A2(n_353),
.B1(n_330),
.B2(n_351),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_380),
.B1(n_371),
.B2(n_373),
.Y(n_386)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_369),
.A2(n_350),
.B(n_325),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_384),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_343),
.B1(n_305),
.B2(n_304),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_370),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_383),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_365),
.B(n_298),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_387),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_375),
.A2(n_284),
.B1(n_362),
.B2(n_363),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_316),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_390),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_361),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_376),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_316),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_392),
.A2(n_236),
.B(n_255),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_385),
.A2(n_384),
.B(n_378),
.Y(n_396)
);

OAI211xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_397),
.B(n_399),
.C(n_400),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_383),
.B(n_376),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_398),
.A2(n_381),
.B(n_316),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_391),
.A2(n_381),
.B(n_364),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_395),
.A2(n_391),
.B1(n_393),
.B2(n_390),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_404),
.Y(n_405)
);

OA21x2_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_398),
.B(n_221),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_394),
.A2(n_285),
.B1(n_244),
.B2(n_196),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_244),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_405),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_403),
.Y(n_409)
);


endmodule