module fake_ariane_352_n_1797 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1797);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1797;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_74),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_22),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_107),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_29),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_42),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_33),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_76),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_61),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_96),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_35),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_50),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_25),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_25),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_94),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_37),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_164),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_45),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_86),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_72),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_144),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_137),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_45),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_100),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_51),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_33),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_21),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_69),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_114),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_27),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_51),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_37),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_80),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_29),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_58),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_120),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_145),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_53),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_62),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_157),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_18),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_85),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_98),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_106),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_49),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_160),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_151),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_46),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_81),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_119),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_112),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_39),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_116),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_6),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_89),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_73),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_78),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_104),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_93),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_101),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_91),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_2),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_141),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_161),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_87),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_121),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_47),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_102),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_31),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_131),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_22),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_139),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_39),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_64),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_136),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_152),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_48),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_12),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_13),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_88),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_15),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_7),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_49),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_105),
.Y(n_321)
);

BUFx8_ASAP7_75t_SL g322 ( 
.A(n_5),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_32),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_35),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_190),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_190),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_267),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_190),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_239),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_171),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_175),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_176),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_190),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_190),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_216),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_327),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_254),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_254),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_239),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_260),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_260),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_254),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_198),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_169),
.B(n_1),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_170),
.B(n_1),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_295),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_199),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_203),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_191),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_177),
.B(n_9),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_210),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_213),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_214),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_319),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_183),
.B(n_9),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_174),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_224),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_203),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_216),
.B(n_10),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_218),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_186),
.B(n_10),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_226),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_191),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_187),
.B(n_13),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_268),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_192),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_218),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_227),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_276),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_276),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_228),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_268),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_193),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_229),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_289),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_167),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_235),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_195),
.B(n_14),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_250),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_256),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_200),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_261),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_206),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_232),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_237),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_238),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_216),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_243),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_271),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_332),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_336),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_348),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_395),
.B(n_286),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_167),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_335),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_349),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_365),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_350),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_377),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_350),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_338),
.B(n_274),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_380),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_396),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_360),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_347),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_R g444 ( 
.A(n_339),
.B(n_192),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_344),
.B(n_345),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_374),
.B(n_286),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_360),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_362),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_387),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

BUFx8_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_185),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_353),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_372),
.B(n_196),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_389),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_390),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_207),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_385),
.B(n_185),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_333),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_395),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_356),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_357),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_208),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_361),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_361),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_R g478 ( 
.A(n_354),
.B(n_320),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_363),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_368),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_368),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_362),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_375),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_286),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_484),
.B(n_364),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_484),
.B(n_369),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_448),
.B(n_370),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_434),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_450),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_444),
.A2(n_399),
.B1(n_382),
.B2(n_388),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_448),
.B(n_371),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_450),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_334),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_448),
.B(n_376),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_391),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_478),
.A2(n_402),
.B1(n_394),
.B2(n_397),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_460),
.B(n_449),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_419),
.A2(n_373),
.B1(n_359),
.B2(n_381),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_455),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_430),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_458),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_466),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_400),
.B1(n_406),
.B2(n_342),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_425),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_392),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_419),
.B(n_408),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_455),
.B(n_217),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_437),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_467),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_R g529 ( 
.A(n_452),
.B(n_393),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_458),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_449),
.B(n_358),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_449),
.B(n_384),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_482),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_414),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_419),
.A2(n_367),
.B1(n_381),
.B2(n_398),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_419),
.B(n_367),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_426),
.B(n_329),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_466),
.B(n_401),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_457),
.B(n_230),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_220),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_419),
.A2(n_245),
.B1(n_252),
.B2(n_258),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_457),
.B(n_401),
.Y(n_552)
);

INVx8_ASAP7_75t_L g553 ( 
.A(n_424),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_418),
.B(n_403),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_403),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_457),
.B(n_404),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_438),
.B(n_233),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_435),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_469),
.B(n_404),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_456),
.B(n_405),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_441),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_456),
.B(n_405),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_464),
.B(n_236),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_473),
.B(n_166),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_441),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_428),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_407),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_435),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_445),
.B(n_407),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

BUFx8_ASAP7_75t_SL g576 ( 
.A(n_454),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_447),
.B(n_409),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_422),
.B(n_246),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_461),
.B(n_409),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_462),
.B(n_320),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_483),
.A2(n_303),
.B1(n_328),
.B2(n_291),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_422),
.B(n_166),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_451),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_463),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_465),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_475),
.B(n_324),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_465),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_470),
.B(n_240),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_422),
.B(n_251),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_471),
.A2(n_281),
.B1(n_301),
.B2(n_278),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_479),
.B(n_375),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_479),
.B(n_379),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_479),
.B(n_379),
.Y(n_600)
);

BUFx4f_ASAP7_75t_L g601 ( 
.A(n_422),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_412),
.B(n_296),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_479),
.B(n_257),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_472),
.B(n_181),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_483),
.B(n_263),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_422),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_422),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_474),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_412),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_433),
.B(n_253),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_474),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_477),
.B(n_269),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_443),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_443),
.A2(n_272),
.B1(n_290),
.B2(n_311),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_446),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_446),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_433),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_433),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_433),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_459),
.A2(n_314),
.B1(n_292),
.B2(n_285),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_433),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_433),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_459),
.B(n_275),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_480),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_436),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_481),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_436),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_481),
.B(n_181),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_436),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_555),
.B(n_182),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_555),
.B(n_182),
.Y(n_635)
);

AND2x6_ASAP7_75t_SL g636 ( 
.A(n_572),
.B(n_270),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_495),
.A2(n_209),
.B1(n_315),
.B2(n_189),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_495),
.A2(n_209),
.B1(n_315),
.B2(n_189),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_531),
.B(n_325),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_498),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_508),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_524),
.B(n_296),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_505),
.B(n_184),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_543),
.B(n_284),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_505),
.B(n_184),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_194),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_533),
.B(n_534),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_533),
.B(n_194),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_534),
.B(n_248),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_248),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_541),
.B(n_323),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_538),
.B(n_323),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_547),
.B(n_298),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_490),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_487),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_489),
.B(n_305),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_313),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_574),
.B(n_316),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_510),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_496),
.B(n_220),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_487),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_538),
.A2(n_277),
.B1(n_326),
.B2(n_283),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_487),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_535),
.B(n_296),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_574),
.B(n_317),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_560),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_503),
.B(n_318),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_506),
.A2(n_287),
.B1(n_293),
.B2(n_302),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_510),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_506),
.A2(n_304),
.B1(n_309),
.B2(n_308),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_578),
.B(n_172),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_500),
.B(n_436),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_521),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_526),
.B(n_279),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_620),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_578),
.B(n_173),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_576),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_489),
.B(n_299),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_520),
.B(n_494),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_612),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_551),
.A2(n_179),
.B1(n_307),
.B2(n_306),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_553),
.B(n_279),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_499),
.B(n_299),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_521),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_501),
.B(n_507),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_612),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_491),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_530),
.B(n_178),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_502),
.B(n_180),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_532),
.B(n_197),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_532),
.B(n_202),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_499),
.A2(n_244),
.B1(n_204),
.B2(n_205),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_560),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_554),
.B(n_211),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_560),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_514),
.B(n_212),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_491),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_509),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_513),
.B(n_215),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_554),
.B(n_221),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_485),
.B(n_14),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_501),
.B(n_507),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_485),
.B(n_15),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_603),
.A2(n_300),
.B1(n_225),
.B2(n_234),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_486),
.A2(n_259),
.B1(n_223),
.B2(n_241),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_513),
.B(n_442),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_516),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_511),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_540),
.B(n_442),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_497),
.B(n_442),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_488),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_497),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_512),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_613),
.A2(n_442),
.B(n_440),
.C(n_436),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_552),
.B(n_273),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_556),
.B(n_265),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_588),
.A2(n_255),
.B1(n_242),
.B2(n_247),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_569),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_618),
.B(n_282),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_486),
.B(n_522),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_618),
.B(n_294),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_512),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_492),
.B(n_442),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_504),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_540),
.B(n_442),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_606),
.B(n_297),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_492),
.B(n_440),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_440),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_526),
.B(n_440),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_522),
.B(n_17),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_515),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_572),
.B(n_19),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_515),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_504),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_606),
.B(n_280),
.Y(n_738)
);

NAND2x1_ASAP7_75t_L g739 ( 
.A(n_621),
.B(n_440),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_551),
.B(n_264),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_557),
.B(n_440),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_558),
.B(n_19),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_518),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_558),
.B(n_20),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_582),
.B(n_20),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_519),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_262),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_525),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_557),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_504),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_593),
.B(n_249),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_570),
.B(n_436),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_528),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_539),
.A2(n_587),
.B1(n_545),
.B2(n_544),
.Y(n_754)
);

BUFx5_ASAP7_75t_L g755 ( 
.A(n_620),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_597),
.B(n_321),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_564),
.B(n_23),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_536),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_570),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_619),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_564),
.B(n_24),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_542),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_582),
.B(n_24),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_604),
.B(n_26),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_550),
.B(n_28),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_559),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_575),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_553),
.B(n_572),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_546),
.A2(n_321),
.B1(n_231),
.B2(n_222),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_549),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_575),
.B(n_321),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_581),
.B(n_28),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_585),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_550),
.B(n_30),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_550),
.B(n_610),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_550),
.B(n_562),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_585),
.B(n_321),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_550),
.B(n_30),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_616),
.A2(n_231),
.B1(n_222),
.B2(n_219),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_591),
.B(n_231),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_568),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_591),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_605),
.B(n_32),
.Y(n_783)
);

BUFx4f_ASAP7_75t_L g784 ( 
.A(n_553),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_596),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_548),
.B(n_34),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_571),
.B(n_34),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_548),
.B(n_38),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_616),
.A2(n_231),
.B1(n_222),
.B2(n_219),
.C(n_201),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_517),
.B(n_577),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_580),
.B(n_38),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_589),
.B(n_41),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_581),
.B(n_231),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_527),
.B(n_222),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_592),
.B(n_41),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_SL g796 ( 
.A(n_596),
.B(n_566),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_594),
.B(n_42),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_602),
.B(n_46),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_609),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_48),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_583),
.A2(n_222),
.B1(n_219),
.B2(n_201),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_649),
.A2(n_561),
.B(n_563),
.C(n_567),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_733),
.A2(n_613),
.B(n_625),
.C(n_584),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_640),
.B(n_628),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_671),
.A2(n_672),
.B1(n_635),
.B2(n_634),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_640),
.B(n_617),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_701),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_654),
.A2(n_632),
.B(n_600),
.C(n_599),
.Y(n_808)
);

AO21x1_ASAP7_75t_L g809 ( 
.A1(n_786),
.A2(n_625),
.B(n_611),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_733),
.A2(n_622),
.B(n_627),
.C(n_630),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_581),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_723),
.B(n_559),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_790),
.A2(n_623),
.B(n_601),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_790),
.A2(n_601),
.B(n_586),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_688),
.B(n_529),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_L g817 ( 
.A1(n_654),
.A2(n_579),
.B(n_595),
.C(n_611),
.Y(n_817)
);

NAND2x1_ASAP7_75t_L g818 ( 
.A(n_796),
.B(n_624),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_678),
.B(n_608),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_742),
.A2(n_744),
.B(n_788),
.C(n_786),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_717),
.A2(n_565),
.B(n_598),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_653),
.A2(n_624),
.B(n_621),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_746),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_653),
.A2(n_565),
.B(n_631),
.Y(n_825)
);

NOR2x1_ASAP7_75t_L g826 ( 
.A(n_680),
.B(n_579),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_672),
.B(n_633),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_664),
.A2(n_629),
.B1(n_607),
.B2(n_608),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_741),
.A2(n_595),
.B(n_608),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_710),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_779),
.A2(n_626),
.B1(n_614),
.B2(n_504),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_650),
.B(n_626),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_741),
.A2(n_608),
.B(n_573),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_752),
.A2(n_573),
.B(n_523),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_698),
.B(n_614),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_651),
.A2(n_52),
.B(n_54),
.C(n_573),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_673),
.A2(n_573),
.B1(n_523),
.B2(n_219),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_723),
.A2(n_523),
.B1(n_219),
.B2(n_201),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_753),
.Y(n_840)
);

OAI321xp33_ASAP7_75t_L g841 ( 
.A1(n_742),
.A2(n_201),
.A3(n_188),
.B1(n_168),
.B2(n_523),
.C(n_52),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_752),
.A2(n_201),
.B(n_188),
.Y(n_842)
);

OAI321xp33_ASAP7_75t_L g843 ( 
.A1(n_744),
.A2(n_188),
.A3(n_168),
.B1(n_54),
.B2(n_63),
.C(n_68),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_644),
.A2(n_188),
.B1(n_168),
.B2(n_79),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_675),
.A2(n_188),
.B(n_168),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_788),
.A2(n_168),
.B(n_57),
.C(n_90),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_783),
.A2(n_55),
.B(n_110),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_696),
.B(n_117),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_675),
.A2(n_124),
.B(n_125),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_704),
.B(n_129),
.C(n_133),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_705),
.B(n_140),
.Y(n_851)
);

NOR2x1_ASAP7_75t_L g852 ( 
.A(n_685),
.B(n_143),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_657),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_678),
.B(n_147),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_784),
.B(n_149),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_690),
.A2(n_150),
.B(n_155),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_696),
.B(n_158),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_661),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_784),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_676),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_685),
.B(n_768),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_762),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_770),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_678),
.B(n_755),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_687),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_781),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_641),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_682),
.A2(n_776),
.B(n_777),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_700),
.A2(n_725),
.B(n_736),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_715),
.A2(n_767),
.B(n_734),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_716),
.A2(n_785),
.B(n_759),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_749),
.A2(n_782),
.B(n_773),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_682),
.A2(n_713),
.B(n_754),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_647),
.B(n_681),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_681),
.B(n_686),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_704),
.A2(n_706),
.B(n_783),
.C(n_658),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_739),
.A2(n_694),
.B(n_691),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_706),
.A2(n_658),
.B(n_791),
.C(n_795),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_693),
.A2(n_728),
.B(n_709),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_678),
.B(n_755),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_709),
.A2(n_712),
.B(n_728),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_686),
.B(n_799),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_712),
.A2(n_648),
.B(n_764),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_678),
.B(n_755),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_791),
.A2(n_795),
.B(n_637),
.C(n_638),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_768),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_768),
.Y(n_887)
);

AO21x1_ASAP7_75t_L g888 ( 
.A1(n_765),
.A2(n_778),
.B(n_774),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_766),
.A2(n_652),
.B(n_719),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_642),
.B(n_643),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_683),
.B(n_689),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_766),
.A2(n_718),
.B(n_668),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_794),
.Y(n_893)
);

BUFx4f_ASAP7_75t_L g894 ( 
.A(n_685),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_731),
.B(n_726),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_771),
.A2(n_777),
.B(n_780),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_787),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_730),
.B(n_656),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_727),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_663),
.A2(n_665),
.B(n_722),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_666),
.B(n_656),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_678),
.B(n_755),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_670),
.B(n_639),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_645),
.B(n_697),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_792),
.A2(n_797),
.B(n_800),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_703),
.B(n_760),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_721),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_760),
.Y(n_908)
);

CKINVDCx10_ASAP7_75t_R g909 ( 
.A(n_758),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_724),
.A2(n_679),
.B(n_674),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_702),
.A2(n_775),
.B(n_738),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_747),
.B(n_751),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_660),
.B(n_667),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_771),
.A2(n_780),
.B(n_756),
.Y(n_914)
);

NOR2x1_ASAP7_75t_L g915 ( 
.A(n_793),
.B(n_735),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_745),
.B(n_763),
.C(n_646),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_745),
.B(n_763),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_793),
.B(n_772),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_793),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_729),
.B(n_662),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_727),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_798),
.A2(n_655),
.B(n_659),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_727),
.A2(n_737),
.B(n_750),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_662),
.B(n_714),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_720),
.B(n_677),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_727),
.A2(n_737),
.B(n_750),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_757),
.B(n_761),
.C(n_699),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_677),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_657),
.B(n_737),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_801),
.A2(n_740),
.B(n_692),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_695),
.A2(n_708),
.B(n_684),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_737),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_636),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_657),
.Y(n_934)
);

NOR2x1_ASAP7_75t_L g935 ( 
.A(n_657),
.B(n_750),
.Y(n_935)
);

OR2x2_ASAP7_75t_SL g936 ( 
.A(n_707),
.B(n_779),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_750),
.A2(n_769),
.B1(n_789),
.B2(n_732),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_732),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_755),
.A2(n_507),
.B(n_501),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_755),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_758),
.B(n_508),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_758),
.A2(n_348),
.B1(n_349),
.B2(n_336),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_649),
.A2(n_671),
.B1(n_672),
.B2(n_634),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_649),
.B(n_493),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_640),
.B(n_649),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_649),
.B(n_493),
.Y(n_949)
);

AOI21xp33_ASAP7_75t_L g950 ( 
.A1(n_681),
.A2(n_529),
.B(n_686),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_649),
.B(n_493),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_796),
.A2(n_675),
.B(n_682),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_710),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_640),
.B(n_649),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_669),
.B(n_698),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_701),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_649),
.B(n_493),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_649),
.B(n_678),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_649),
.B(n_671),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_796),
.A2(n_675),
.B(n_682),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_669),
.B(n_698),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_649),
.B(n_671),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_649),
.B(n_493),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_701),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_710),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_640),
.B(n_649),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_701),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_649),
.B(n_493),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_649),
.A2(n_671),
.B1(n_672),
.B2(n_634),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_701),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_727),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_758),
.B(n_508),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_640),
.B(n_649),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_649),
.B(n_671),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_723),
.A2(n_495),
.B1(n_733),
.B2(n_706),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_649),
.B(n_493),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_758),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_688),
.B(n_531),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_649),
.B(n_493),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_796),
.A2(n_675),
.B(n_682),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_654),
.A2(n_419),
.B1(n_551),
.B2(n_664),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_649),
.A2(n_671),
.B1(n_672),
.B2(n_634),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_649),
.A2(n_790),
.B(n_653),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_876),
.A2(n_878),
.B(n_941),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_858),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_960),
.A2(n_947),
.B(n_942),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_853),
.Y(n_993)
);

OAI22x1_ASAP7_75t_L g994 ( 
.A1(n_979),
.A2(n_918),
.B1(n_906),
.B2(n_915),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_853),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_948),
.B(n_956),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_867),
.Y(n_997)
);

AND3x2_ASAP7_75t_L g998 ( 
.A(n_925),
.B(n_893),
.C(n_931),
.Y(n_998)
);

AOI221xp5_ASAP7_75t_SL g999 ( 
.A1(n_885),
.A2(n_820),
.B1(n_803),
.B2(n_964),
.C(n_961),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_984),
.A2(n_888),
.B(n_873),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_860),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_954),
.A2(n_967),
.B(n_955),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_969),
.A2(n_988),
.B(n_986),
.Y(n_1003)
);

AO31x2_ASAP7_75t_L g1004 ( 
.A1(n_809),
.A2(n_810),
.A3(n_896),
.B(n_883),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_909),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_900),
.A2(n_880),
.B(n_864),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_864),
.A2(n_884),
.B(n_880),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_917),
.A2(n_875),
.B1(n_961),
.B2(n_978),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_879),
.A2(n_914),
.B(n_817),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_964),
.A2(n_978),
.B(n_956),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_831),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_817),
.A2(n_845),
.B(n_892),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_948),
.A2(n_977),
.B(n_970),
.C(n_950),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_865),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_812),
.B(n_945),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_877),
.A2(n_819),
.B(n_911),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_821),
.A2(n_902),
.B(n_884),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_902),
.A2(n_926),
.B(n_923),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_819),
.A2(n_889),
.B(n_910),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_970),
.A2(n_977),
.B(n_874),
.C(n_841),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_946),
.A2(n_972),
.B1(n_965),
.B2(n_959),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_881),
.A2(n_834),
.B(n_835),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_814),
.A2(n_849),
.B(n_854),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_812),
.B(n_973),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_949),
.A2(n_983),
.B(n_980),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_951),
.B(n_816),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_807),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_912),
.B(n_906),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_912),
.B(n_882),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_903),
.B(n_893),
.Y(n_1030)
);

AOI221x1_ASAP7_75t_L g1031 ( 
.A1(n_847),
.A2(n_927),
.B1(n_916),
.B2(n_844),
.C(n_805),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_987),
.A2(n_930),
.B(n_854),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_842),
.A2(n_830),
.B(n_905),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_813),
.A2(n_828),
.B(n_833),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_982),
.B(n_913),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_802),
.A2(n_822),
.B(n_895),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_985),
.A2(n_897),
.B1(n_974),
.B2(n_862),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_908),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_815),
.B(n_823),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_808),
.A2(n_940),
.B(n_922),
.Y(n_1040)
);

AO21x2_ASAP7_75t_L g1041 ( 
.A1(n_927),
.A2(n_825),
.B(n_839),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_944),
.B(n_908),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_829),
.A2(n_818),
.B(n_870),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_953),
.B(n_924),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_859),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_869),
.A2(n_871),
.B(n_872),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_L g1047 ( 
.A(n_943),
.B(n_976),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_853),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_929),
.A2(n_935),
.B(n_898),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_981),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_824),
.Y(n_1051)
);

CKINVDCx8_ASAP7_75t_R g1052 ( 
.A(n_932),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_827),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_929),
.A2(n_856),
.B(n_975),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_899),
.A2(n_975),
.B(n_921),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_899),
.A2(n_921),
.B(n_934),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_SL g1057 ( 
.A(n_855),
.B(n_853),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_886),
.B(n_938),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_838),
.A2(n_843),
.B(n_901),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_985),
.A2(n_904),
.B(n_937),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_840),
.B(n_971),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_837),
.A2(n_850),
.B(n_806),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_804),
.A2(n_852),
.B(n_832),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_863),
.B(n_866),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_891),
.A2(n_966),
.B(n_958),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_920),
.B(n_939),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_836),
.B(n_919),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_851),
.A2(n_832),
.B(n_861),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_957),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_846),
.A2(n_848),
.B(n_857),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_968),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_957),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_894),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_848),
.B(n_857),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_890),
.A2(n_938),
.B(n_907),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_963),
.B(n_928),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_963),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_936),
.A2(n_886),
.B(n_811),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_938),
.A2(n_826),
.A3(n_887),
.B(n_894),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_811),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_933),
.A2(n_917),
.B1(n_878),
.B2(n_979),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_831),
.B(n_553),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_876),
.A2(n_649),
.B(n_878),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_909),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_952),
.A2(n_984),
.B(n_962),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_875),
.A2(n_874),
.B(n_917),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_807),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_888),
.A2(n_809),
.A3(n_820),
.B(n_876),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_807),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_876),
.B(n_878),
.C(n_979),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_816),
.B(n_450),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_867),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_876),
.A2(n_649),
.B(n_878),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_979),
.A2(n_820),
.B(n_876),
.C(n_878),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_820),
.B(n_876),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_SL g1107 ( 
.A1(n_820),
.A2(n_876),
.B(n_878),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_979),
.A2(n_820),
.B(n_876),
.C(n_878),
.Y(n_1108)
);

AOI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_875),
.A2(n_529),
.B(n_430),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_979),
.A2(n_820),
.B(n_876),
.C(n_878),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_917),
.A2(n_875),
.B(n_874),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_868),
.A2(n_962),
.B(n_952),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_868),
.A2(n_984),
.B(n_962),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_952),
.A2(n_984),
.B(n_962),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_816),
.B(n_569),
.Y(n_1115)
);

AND2x2_ASAP7_75t_SL g1116 ( 
.A(n_894),
.B(n_875),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_807),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_948),
.B(n_956),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_831),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_858),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_932),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_979),
.A2(n_820),
.B(n_876),
.C(n_878),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_908),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_868),
.A2(n_984),
.B(n_962),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_948),
.B(n_956),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_875),
.A2(n_529),
.B(n_430),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_960),
.A2(n_649),
.B(n_941),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_868),
.A2(n_984),
.B(n_962),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_952),
.A2(n_984),
.B(n_962),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_858),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_876),
.A2(n_649),
.B(n_878),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_948),
.B(n_956),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_SL g1138 ( 
.A1(n_979),
.A2(n_910),
.B(n_881),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_948),
.B(n_956),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_979),
.A2(n_820),
.B(n_876),
.C(n_878),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_888),
.A2(n_809),
.A3(n_820),
.B(n_876),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_996),
.B(n_1120),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_993),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1070),
.A2(n_1024),
.B(n_1015),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1129),
.B(n_1137),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1038),
.B(n_1126),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1038),
.B(n_1126),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1074),
.A2(n_1028),
.B1(n_1081),
.B2(n_1139),
.Y(n_1148)
);

BUFx4f_ASAP7_75t_L g1149 ( 
.A(n_1082),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_997),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_993),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1121),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1015),
.A2(n_1024),
.B(n_1025),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_993),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1005),
.Y(n_1155)
);

BUFx2_ASAP7_75t_SL g1156 ( 
.A(n_1052),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1099),
.B(n_1035),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_SL g1158 ( 
.A(n_1084),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1021),
.A2(n_1102),
.B(n_1083),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1013),
.B(n_1029),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1073),
.B(n_1123),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1116),
.A2(n_1097),
.B1(n_994),
.B2(n_1042),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1101),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_1097),
.A2(n_1010),
.B1(n_1136),
.B2(n_1104),
.C1(n_1008),
.C2(n_1108),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1072),
.B(n_1115),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1103),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1116),
.A2(n_999),
.B1(n_1109),
.B2(n_1130),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1030),
.B(n_998),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1027),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_SL g1171 ( 
.A1(n_1104),
.A2(n_990),
.B(n_1037),
.C(n_1117),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1051),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1123),
.B(n_1121),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1050),
.B(n_1011),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_995),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1082),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1053),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1103),
.A2(n_1125),
.B1(n_1110),
.B2(n_1108),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1110),
.A2(n_1140),
.B(n_1020),
.C(n_1138),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_1005),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1044),
.B(n_1072),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1079),
.B(n_1082),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1140),
.B(n_1020),
.C(n_1031),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1059),
.A2(n_1060),
.B(n_1066),
.C(n_1062),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1086),
.B(n_998),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1039),
.A2(n_1064),
.B1(n_1061),
.B2(n_1087),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1071),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1095),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1001),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1071),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1014),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1079),
.B(n_1069),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1045),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1076),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1062),
.A2(n_1017),
.B(n_1055),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1002),
.A2(n_1003),
.B(n_1118),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1077),
.B(n_1122),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1067),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1080),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1045),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_L g1201 ( 
.A(n_992),
.B(n_1040),
.C(n_1088),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1080),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1066),
.A2(n_1065),
.B(n_1075),
.C(n_1063),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_995),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1032),
.A2(n_1119),
.B(n_1132),
.C(n_1124),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1058),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1135),
.B(n_1078),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1036),
.A2(n_1131),
.B(n_1127),
.C(n_1100),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1079),
.B(n_1047),
.Y(n_1209)
);

BUFx4_ASAP7_75t_SL g1210 ( 
.A(n_1057),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1089),
.A2(n_1034),
.B1(n_1058),
.B2(n_1048),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1068),
.A2(n_1041),
.B1(n_1063),
.B2(n_1048),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_1023),
.B(n_1006),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1093),
.B(n_1141),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1041),
.A2(n_1111),
.B(n_1046),
.C(n_1093),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1049),
.B(n_1056),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1007),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1093),
.Y(n_1218)
);

BUFx5_ASAP7_75t_L g1219 ( 
.A(n_1085),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1009),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1111),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1017),
.A2(n_1023),
.B1(n_1054),
.B2(n_1033),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1141),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1141),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1018),
.B(n_1033),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1004),
.B(n_1009),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1004),
.B(n_1000),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1018),
.B(n_989),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1004),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1090),
.B(n_1105),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1114),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1019),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1022),
.A2(n_1012),
.B(n_1106),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1113),
.B(n_1128),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1134),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1091),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1016),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1133),
.A2(n_1092),
.B(n_1094),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1112),
.C(n_1133),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1012),
.A2(n_1070),
.B(n_1024),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1121),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_996),
.B(n_1120),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_997),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1005),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1082),
.Y(n_1245)
);

CKINVDCx8_ASAP7_75t_R g1246 ( 
.A(n_1005),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1038),
.B(n_903),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1011),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_996),
.B(n_1120),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1070),
.A2(n_1024),
.B(n_1015),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1027),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_996),
.B(n_1120),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1074),
.A2(n_875),
.B1(n_588),
.B2(n_979),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1015),
.A2(n_1024),
.B(n_1104),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1011),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_997),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1082),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1121),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_996),
.B(n_1120),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_991),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1005),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1073),
.B(n_886),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1073),
.B(n_886),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1074),
.B(n_1028),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_990),
.A2(n_1107),
.B(n_1083),
.C(n_1102),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1038),
.B(n_903),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1038),
.B(n_903),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1027),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1070),
.A2(n_1024),
.B(n_1015),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1074),
.A2(n_360),
.B1(n_362),
.B2(n_350),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1073),
.B(n_886),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1027),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1074),
.A2(n_979),
.B1(n_1028),
.B2(n_878),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1070),
.A2(n_1024),
.B(n_1015),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1073),
.B(n_886),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1070),
.A2(n_1024),
.B(n_1015),
.Y(n_1277)
);

BUFx5_ASAP7_75t_L g1278 ( 
.A(n_1116),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_SL g1279 ( 
.A1(n_1104),
.A2(n_990),
.B(n_1081),
.C(n_1024),
.Y(n_1279)
);

OAI31xp33_ASAP7_75t_L g1280 ( 
.A1(n_1081),
.A2(n_820),
.A3(n_1028),
.B(n_878),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1146),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1169),
.A2(n_1185),
.B1(n_1183),
.B2(n_1157),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1248),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1185),
.A2(n_1183),
.B1(n_1280),
.B2(n_1161),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1233),
.A2(n_1213),
.B(n_1205),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1178),
.A2(n_1274),
.B1(n_1161),
.B2(n_1160),
.Y(n_1286)
);

INVxp33_ASAP7_75t_L g1287 ( 
.A(n_1257),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1196),
.A2(n_1240),
.B(n_1201),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1175),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1196),
.A2(n_1239),
.B(n_1215),
.Y(n_1290)
);

BUFx5_ASAP7_75t_L g1291 ( 
.A(n_1216),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1254),
.A2(n_1148),
.B1(n_1163),
.B2(n_1253),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1246),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1155),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1201),
.A2(n_1184),
.B(n_1144),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1259),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1170),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1214),
.B(n_1147),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1190),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1237),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1182),
.B(n_1209),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1172),
.Y(n_1302)
);

INVxp67_ASAP7_75t_SL g1303 ( 
.A(n_1186),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1247),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1251),
.A2(n_1270),
.B(n_1277),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1173),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1177),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1156),
.A2(n_1142),
.B1(n_1260),
.B2(n_1145),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1180),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1188),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1244),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1218),
.B(n_1223),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1280),
.A2(n_1274),
.B1(n_1160),
.B2(n_1271),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1212),
.A2(n_1203),
.B(n_1207),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1252),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1269),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1262),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1229),
.A2(n_1167),
.B1(n_1159),
.B2(n_1192),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1178),
.A2(n_1186),
.B1(n_1275),
.B2(n_1149),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1153),
.A2(n_1222),
.B(n_1234),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1174),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1209),
.B(n_1182),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1142),
.B(n_1145),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1165),
.A2(n_1179),
.B(n_1168),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1273),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1211),
.A2(n_1255),
.B(n_1234),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1197),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1189),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1191),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1195),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1258),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1158),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1261),
.Y(n_1333)
);

AOI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1211),
.A2(n_1225),
.B(n_1231),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1242),
.B(n_1250),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1200),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1230),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1158),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1149),
.A2(n_1194),
.B1(n_1258),
.B2(n_1278),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1267),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1268),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1225),
.A2(n_1235),
.B(n_1228),
.Y(n_1342)
);

CKINVDCx16_ASAP7_75t_R g1343 ( 
.A(n_1173),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1230),
.Y(n_1344)
);

INVx8_ASAP7_75t_L g1345 ( 
.A(n_1263),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1165),
.A2(n_1207),
.B1(n_1253),
.B2(n_1242),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1250),
.B(n_1260),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1278),
.A2(n_1198),
.B1(n_1166),
.B2(n_1245),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1181),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1224),
.B(n_1227),
.Y(n_1350)
);

CKINVDCx11_ASAP7_75t_R g1351 ( 
.A(n_1150),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1224),
.B(n_1279),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1265),
.B(n_1278),
.Y(n_1353)
);

CKINVDCx14_ASAP7_75t_R g1354 ( 
.A(n_1249),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1150),
.A2(n_1243),
.B1(n_1164),
.B2(n_1221),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1278),
.A2(n_1243),
.B1(n_1164),
.B2(n_1199),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1256),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1152),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1187),
.A2(n_1193),
.B1(n_1245),
.B2(n_1266),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1278),
.B(n_1143),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1176),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1143),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1204),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1238),
.A2(n_1226),
.B(n_1208),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1151),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1241),
.A2(n_1199),
.B1(n_1202),
.B2(n_1162),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1162),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1219),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1206),
.A2(n_1276),
.B1(n_1272),
.B2(n_1263),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1264),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1154),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1264),
.B(n_1276),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1272),
.B(n_1171),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1236),
.Y(n_1376)
);

BUFx2_ASAP7_75t_R g1377 ( 
.A(n_1210),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1217),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1220),
.B2(n_1219),
.Y(n_1379)
);

BUFx8_ASAP7_75t_SL g1380 ( 
.A(n_1232),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1220),
.A2(n_950),
.B1(n_336),
.B2(n_349),
.Y(n_1381)
);

BUFx8_ASAP7_75t_SL g1382 ( 
.A(n_1180),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1170),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1170),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1237),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1163),
.A2(n_643),
.B1(n_666),
.B2(n_1074),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1170),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1180),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1233),
.A2(n_1213),
.B(n_1205),
.Y(n_1389)
);

INVx4_ASAP7_75t_SL g1390 ( 
.A(n_1229),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1237),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1170),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1175),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1148),
.A2(n_1074),
.B1(n_1254),
.B2(n_979),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1170),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1213),
.A2(n_1233),
.B(n_1003),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1175),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1396),
.A2(n_1389),
.B(n_1285),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1376),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1337),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1298),
.B(n_1350),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1323),
.B(n_1321),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1298),
.B(n_1281),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1303),
.B(n_1346),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1286),
.B(n_1284),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1337),
.B(n_1344),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1328),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1329),
.Y(n_1408)
);

AOI21xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1394),
.A2(n_1292),
.B(n_1386),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1396),
.A2(n_1389),
.B(n_1285),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1299),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1335),
.B(n_1347),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1308),
.B(n_1319),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1290),
.A2(n_1330),
.B(n_1365),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1380),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1352),
.A2(n_1334),
.B(n_1326),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1312),
.B(n_1304),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1312),
.B(n_1297),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1378),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1302),
.B(n_1307),
.Y(n_1422)
);

BUFx4f_ASAP7_75t_SL g1423 ( 
.A(n_1388),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1288),
.Y(n_1425)
);

INVx4_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1316),
.B(n_1325),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1383),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1290),
.A2(n_1330),
.B(n_1365),
.Y(n_1429)
);

OAI21xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1313),
.A2(n_1353),
.B(n_1318),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1324),
.A2(n_1375),
.B(n_1295),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1295),
.A2(n_1359),
.B(n_1305),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1288),
.A2(n_1295),
.B(n_1320),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1288),
.A2(n_1320),
.B(n_1305),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1384),
.Y(n_1435)
);

NAND2x1_ASAP7_75t_L g1436 ( 
.A(n_1305),
.B(n_1368),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1291),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1368),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1387),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1392),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1361),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1395),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1353),
.B(n_1340),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1370),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1314),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1341),
.B(n_1301),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1314),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1306),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1360),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1355),
.A2(n_1381),
.B(n_1367),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1300),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1349),
.B(n_1300),
.Y(n_1454)
);

NAND2x1_ASAP7_75t_L g1455 ( 
.A(n_1360),
.B(n_1379),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1282),
.A2(n_1287),
.B(n_1391),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1333),
.A2(n_1373),
.B(n_1366),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1385),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1385),
.B(n_1391),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1322),
.B(n_1327),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1287),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1354),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1437),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1401),
.B(n_1362),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1415),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1403),
.B(n_1343),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1415),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1409),
.A2(n_1369),
.B1(n_1339),
.B2(n_1371),
.C(n_1283),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1400),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1457),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1403),
.B(n_1358),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1401),
.B(n_1362),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1409),
.B(n_1351),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1419),
.B(n_1358),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1436),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1419),
.B(n_1283),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1457),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1407),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1405),
.A2(n_1351),
.B1(n_1345),
.B2(n_1374),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1407),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1451),
.B(n_1354),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1433),
.B(n_1364),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1451),
.B(n_1364),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.B(n_1425),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1431),
.B(n_1289),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1408),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1289),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1405),
.A2(n_1345),
.B1(n_1331),
.B2(n_1357),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1289),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1431),
.A2(n_1390),
.B(n_1331),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1452),
.A2(n_1345),
.B1(n_1372),
.B2(n_1357),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1438),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1417),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1415),
.B(n_1397),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1421),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1404),
.B(n_1393),
.Y(n_1498)
);

OAI211xp5_ASAP7_75t_L g1499 ( 
.A1(n_1414),
.A2(n_1452),
.B(n_1404),
.C(n_1432),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1421),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1498),
.B(n_1412),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1498),
.B(n_1439),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1474),
.A2(n_1414),
.B1(n_1458),
.B2(n_1402),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1406),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1479),
.Y(n_1505)
);

OAI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1469),
.A2(n_1463),
.B1(n_1456),
.B2(n_1489),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1499),
.A2(n_1430),
.B1(n_1458),
.B2(n_1463),
.C(n_1454),
.Y(n_1508)
);

OAI21xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1482),
.A2(n_1474),
.B(n_1467),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1469),
.A2(n_1430),
.B1(n_1456),
.B2(n_1460),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1497),
.B(n_1461),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1489),
.B(n_1406),
.Y(n_1512)
);

NAND2x1_ASAP7_75t_L g1513 ( 
.A(n_1464),
.B(n_1400),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1500),
.B(n_1453),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1466),
.A2(n_1434),
.B(n_1398),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1466),
.A2(n_1398),
.B(n_1411),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1500),
.B(n_1499),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1493),
.A2(n_1413),
.B1(n_1454),
.B2(n_1428),
.C(n_1435),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1420),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1492),
.A2(n_1468),
.B1(n_1466),
.B2(n_1445),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1468),
.A2(n_1413),
.B1(n_1428),
.B2(n_1440),
.C(n_1435),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1475),
.B(n_1459),
.C(n_1416),
.D(n_1426),
.Y(n_1522)
);

OAI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1493),
.A2(n_1443),
.B1(n_1440),
.B2(n_1441),
.C(n_1455),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1473),
.B(n_1420),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1471),
.A2(n_1441),
.B1(n_1443),
.B2(n_1427),
.C(n_1424),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1471),
.A2(n_1427),
.B1(n_1424),
.B2(n_1422),
.C(n_1445),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1480),
.A2(n_1416),
.B1(n_1426),
.B2(n_1462),
.Y(n_1527)
);

OAI21xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1482),
.A2(n_1459),
.B(n_1416),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1473),
.B(n_1442),
.Y(n_1529)
);

OAI21xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1482),
.A2(n_1467),
.B(n_1426),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_R g1531 ( 
.A(n_1467),
.B(n_1332),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1486),
.B(n_1450),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1480),
.A2(n_1416),
.B1(n_1426),
.B2(n_1423),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1490),
.B(n_1429),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1477),
.A2(n_1475),
.B1(n_1472),
.B2(n_1486),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1485),
.A2(n_1410),
.B(n_1399),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1490),
.B(n_1484),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1477),
.B(n_1332),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1465),
.B(n_1422),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1465),
.B(n_1448),
.Y(n_1540)
);

NOR3xp33_ASAP7_75t_SL g1541 ( 
.A(n_1495),
.B(n_1293),
.C(n_1338),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1478),
.A2(n_1449),
.B1(n_1447),
.B2(n_1460),
.C(n_1418),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1472),
.B(n_1446),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1490),
.B(n_1429),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1507),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1514),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1534),
.B(n_1545),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1528),
.B(n_1475),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1502),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1517),
.B(n_1491),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1501),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1537),
.B(n_1483),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1476),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1525),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1539),
.B(n_1472),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1504),
.B(n_1483),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1515),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1516),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1491),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1543),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1535),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1519),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1532),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1542),
.B(n_1494),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1516),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_1496),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1508),
.A2(n_1477),
.B1(n_1494),
.B2(n_1429),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1566),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1546),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1562),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1547),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1556),
.B(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1547),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1479),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1548),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1555),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1580),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1562),
.B(n_1338),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1580),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1575),
.B(n_1309),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1550),
.B(n_1481),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1550),
.B(n_1481),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1551),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1538),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1560),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1569),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1570),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1551),
.B(n_1481),
.Y(n_1612)
);

INVx5_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1560),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1568),
.B(n_1518),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1570),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1572),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1574),
.B(n_1450),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1585),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1588),
.B(n_1579),
.C(n_1574),
.D(n_1527),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1588),
.B(n_1576),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1592),
.B(n_1576),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1583),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1613),
.B(n_1561),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1583),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1613),
.B(n_1561),
.Y(n_1628)
);

NAND4xp25_ASAP7_75t_L g1629 ( 
.A(n_1600),
.B(n_1579),
.C(n_1533),
.D(n_1578),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_SL g1631 ( 
.A(n_1586),
.B(n_1578),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1613),
.B(n_1575),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1613),
.B(n_1560),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1568),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1589),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1613),
.B(n_1559),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1581),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1589),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1594),
.B(n_1581),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1591),
.Y(n_1643)
);

OAI31xp33_ASAP7_75t_L g1644 ( 
.A1(n_1616),
.A2(n_1506),
.A3(n_1523),
.B(n_1565),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1611),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1597),
.B(n_1309),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1613),
.B(n_1553),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1591),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1616),
.A2(n_1565),
.B(n_1520),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1619),
.B(n_1567),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_SL g1654 ( 
.A(n_1619),
.B(n_1377),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1596),
.B(n_1573),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_SL g1656 ( 
.A1(n_1607),
.A2(n_1388),
.B(n_1563),
.C(n_1573),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1563),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1605),
.B(n_1552),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1619),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1584),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1590),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1602),
.B(n_1564),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1623),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1635),
.B(n_1618),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1623),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1621),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1621),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1646),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1647),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1586),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1661),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1630),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1626),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1382),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1598),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1636),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1650),
.A2(n_1492),
.B1(n_1510),
.B2(n_1620),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1640),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1647),
.Y(n_1684)
);

INVxp33_ASAP7_75t_L g1685 ( 
.A(n_1622),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1624),
.B(n_1382),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1643),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1632),
.A2(n_1577),
.B(n_1557),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1598),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1606),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1626),
.B(n_1606),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1633),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1631),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1644),
.B(n_1618),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1633),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1599),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1641),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1685),
.B(n_1629),
.C(n_1643),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1667),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1667),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1668),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1662),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1669),
.B(n_1656),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1694),
.B(n_1695),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

OAI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1699),
.A2(n_1631),
.B(n_1628),
.Y(n_1709)
);

AOI322xp5_ASAP7_75t_L g1710 ( 
.A1(n_1682),
.A2(n_1549),
.A3(n_1557),
.B1(n_1577),
.B2(n_1645),
.C1(n_1627),
.C2(n_1653),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1694),
.A2(n_1627),
.B1(n_1625),
.B2(n_1642),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1673),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1648),
.C(n_1662),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1673),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1666),
.B(n_1599),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1696),
.A2(n_1557),
.B1(n_1549),
.B2(n_1653),
.C(n_1642),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1688),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1688),
.A2(n_1652),
.B1(n_1625),
.B2(n_1645),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1549),
.C(n_1638),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1690),
.B(n_1610),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1617),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1677),
.Y(n_1723)
);

OAI322xp33_ASAP7_75t_L g1724 ( 
.A1(n_1678),
.A2(n_1657),
.A3(n_1655),
.B1(n_1648),
.B2(n_1659),
.C1(n_1660),
.C2(n_1651),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1684),
.A2(n_1671),
.B(n_1697),
.C(n_1693),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1702),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1706),
.B(n_1686),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1293),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1701),
.B(n_1689),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1711),
.B(n_1665),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1718),
.A2(n_1638),
.B1(n_1652),
.B2(n_1671),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1718),
.A2(n_1492),
.B1(n_1688),
.B2(n_1692),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1707),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1678),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1703),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1721),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1704),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1708),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1716),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1722),
.B(n_1698),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1725),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1713),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1709),
.B(n_1675),
.Y(n_1744)
);

AOI222xp33_ASAP7_75t_L g1745 ( 
.A1(n_1719),
.A2(n_1687),
.B1(n_1680),
.B2(n_1681),
.C1(n_1677),
.C2(n_1679),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1733),
.B(n_1693),
.Y(n_1746)
);

AO21x1_ASAP7_75t_L g1747 ( 
.A1(n_1736),
.A2(n_1723),
.B(n_1715),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1733),
.B(n_1693),
.Y(n_1748)
);

OAI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1728),
.A2(n_1674),
.B(n_1714),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_SL g1750 ( 
.A(n_1745),
.B(n_1719),
.C(n_1720),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1734),
.A2(n_1731),
.B1(n_1724),
.B2(n_1717),
.C(n_1732),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1728),
.A2(n_1720),
.B(n_1712),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1740),
.A2(n_1735),
.B1(n_1742),
.B2(n_1737),
.C(n_1741),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1730),
.B(n_1698),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1727),
.A2(n_1679),
.B1(n_1680),
.B2(n_1681),
.C(n_1683),
.Y(n_1756)
);

O2A1O1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1743),
.A2(n_1683),
.B(n_1687),
.C(n_1688),
.Y(n_1757)
);

NOR2xp67_ASAP7_75t_L g1758 ( 
.A(n_1752),
.B(n_1743),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1747),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1750),
.A2(n_1738),
.B(n_1736),
.Y(n_1760)
);

AND5x1_ASAP7_75t_L g1761 ( 
.A(n_1751),
.B(n_1744),
.C(n_1710),
.D(n_1693),
.E(n_1697),
.Y(n_1761)
);

NAND4xp75_ASAP7_75t_L g1762 ( 
.A(n_1754),
.B(n_1738),
.C(n_1739),
.D(n_1726),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1749),
.A2(n_1674),
.B1(n_1660),
.B2(n_1628),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1757),
.B(n_1637),
.C(n_1294),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1753),
.B(n_1658),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1755),
.B(n_1633),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1759),
.B(n_1756),
.C(n_1748),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1758),
.B(n_1746),
.Y(n_1768)
);

AOI222xp33_ASAP7_75t_L g1769 ( 
.A1(n_1760),
.A2(n_1764),
.B1(n_1761),
.B2(n_1766),
.C1(n_1763),
.C2(n_1762),
.Y(n_1769)
);

NAND4xp25_ASAP7_75t_SL g1770 ( 
.A(n_1760),
.B(n_1765),
.C(n_1637),
.D(n_1336),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1759),
.A2(n_1294),
.B(n_1633),
.C(n_1655),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1768),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1767),
.Y(n_1773)
);

O2A1O1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1769),
.A2(n_1336),
.B(n_1657),
.C(n_1617),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1770),
.Y(n_1775)
);

AO22x1_ASAP7_75t_L g1776 ( 
.A1(n_1771),
.A2(n_1317),
.B1(n_1311),
.B2(n_1658),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1768),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1777),
.B(n_1531),
.C(n_1296),
.Y(n_1778)
);

NAND4xp75_ASAP7_75t_L g1779 ( 
.A(n_1772),
.B(n_1773),
.C(n_1775),
.D(n_1774),
.Y(n_1779)
);

OAI311xp33_ASAP7_75t_L g1780 ( 
.A1(n_1776),
.A2(n_1614),
.A3(n_1608),
.B1(n_1609),
.C1(n_1593),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1773),
.A2(n_1609),
.B(n_1608),
.Y(n_1781)
);

BUFx2_ASAP7_75t_SL g1782 ( 
.A(n_1777),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1782),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1779),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1781),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1783),
.Y(n_1786)
);

NOR4xp25_ASAP7_75t_L g1787 ( 
.A(n_1786),
.B(n_1784),
.C(n_1785),
.D(n_1780),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1787),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1787),
.Y(n_1789)
);

INVxp33_ASAP7_75t_SL g1790 ( 
.A(n_1788),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1789),
.A2(n_1784),
.B(n_1783),
.Y(n_1791)
);

XNOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1790),
.B(n_1778),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1791),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1792),
.B(n_1317),
.Y(n_1794)
);

AOI222xp33_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1311),
.B1(n_1296),
.B2(n_1552),
.C1(n_1603),
.C2(n_1604),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_R g1796 ( 
.A1(n_1795),
.A2(n_1541),
.B1(n_1607),
.B2(n_1615),
.C(n_1552),
.Y(n_1796)
);

AOI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1399),
.B(n_1410),
.C(n_1612),
.Y(n_1797)
);


endmodule