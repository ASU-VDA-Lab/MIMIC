module fake_jpeg_12834_n_291 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_252;
wire n_251;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_86;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_273;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_26),
.B1(n_19),
.B2(n_38),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_26),
.B1(n_19),
.B2(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_30),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_30),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_20),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_64),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_68),
.B1(n_27),
.B2(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_74),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_28),
.B1(n_18),
.B2(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_28),
.B1(n_18),
.B2(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_36),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_6),
.B(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_84),
.Y(n_140)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_94),
.Y(n_127)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_100),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_96),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_60),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_75),
.B1(n_71),
.B2(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_16),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_33),
.B1(n_1),
.B2(n_4),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_113),
.B1(n_84),
.B2(n_83),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_66),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_16),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_9),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_75),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_117),
.A2(n_123),
.B1(n_78),
.B2(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_90),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_33),
.B(n_71),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_121),
.B(n_134),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_71),
.B(n_33),
.C(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_107),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_132),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_5),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_83),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_9),
.C(n_10),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_89),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_101),
.B1(n_112),
.B2(n_91),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_148),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_132),
.C(n_125),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_81),
.B1(n_101),
.B2(n_103),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_172),
.B1(n_125),
.B2(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_161),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_117),
.B1(n_126),
.B2(n_124),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_97),
.B(n_106),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_155),
.B(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_13),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_97),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_14),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_134),
.B(n_169),
.Y(n_190)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_175),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_130),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_191),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_196),
.B(n_166),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_115),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_168),
.C(n_174),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_128),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_146),
.C(n_158),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_144),
.B1(n_131),
.B2(n_133),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_192),
.B1(n_148),
.B2(n_149),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_199),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_121),
.B(n_137),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_165),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_204),
.B1(n_222),
.B2(n_167),
.Y(n_240)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_149),
.Y(n_208)
);

XOR2x2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_187),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_223),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_147),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_178),
.C(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_180),
.B(n_168),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_217),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_173),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_222),
.B1(n_196),
.B2(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_170),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_204),
.A2(n_172),
.B1(n_179),
.B2(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_203),
.B1(n_209),
.B2(n_207),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_156),
.B(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_202),
.B(n_207),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_198),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_199),
.B1(n_194),
.B2(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_255),
.B1(n_250),
.B2(n_190),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_141),
.B1(n_124),
.B2(n_234),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_246),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_156),
.B(n_223),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_254),
.B(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_158),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_211),
.C(n_212),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_175),
.C(n_126),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_160),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_176),
.C(n_197),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_205),
.B1(n_123),
.B2(n_176),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_264),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_245),
.B1(n_247),
.B2(n_254),
.Y(n_260)
);

NAND4xp25_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.C(n_266),
.D(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_239),
.B1(n_232),
.B2(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_241),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_273),
.B(n_251),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g270 ( 
.A(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_271),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_266),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_279),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_258),
.B1(n_263),
.B2(n_265),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_278),
.B1(n_108),
.B2(n_86),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_10),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_260),
.B1(n_250),
.B2(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_108),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_86),
.C(n_98),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.C(n_98),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_278),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.C(n_282),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_280),
.C(n_11),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_287),
.Y(n_291)
);


endmodule