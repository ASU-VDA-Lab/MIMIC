module fake_jpeg_8242_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_19),
.B1(n_31),
.B2(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_49),
.B1(n_57),
.B2(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_19),
.B1(n_25),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_56),
.B1(n_21),
.B2(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_22),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_15),
.B1(n_29),
.B2(n_17),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_23),
.B1(n_18),
.B2(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_1),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_64),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_14),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_13),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_59),
.C(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_92),
.C(n_21),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_91),
.B(n_1),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_57),
.B1(n_48),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_93),
.B1(n_63),
.B2(n_65),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_57),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_57),
.B(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_74),
.B1(n_68),
.B2(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_66),
.B1(n_62),
.B2(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_108),
.B(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_112),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_77),
.B(n_71),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_39),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_30),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_94),
.B(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_91),
.B1(n_96),
.B2(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_85),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_100),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_91),
.B1(n_84),
.B2(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_80),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_129),
.B(n_110),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_94),
.A3(n_81),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_80),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_101),
.C(n_102),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_1),
.B(n_2),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_138),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_115),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_136),
.C(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_126),
.B1(n_124),
.B2(n_58),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_99),
.B(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_141),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_73),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_125),
.C(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_116),
.B1(n_127),
.B2(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_120),
.C(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_118),
.C(n_130),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_150),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_138),
.B1(n_140),
.B2(n_131),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_153),
.A2(n_52),
.B1(n_6),
.B2(n_8),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_145),
.A2(n_140),
.B(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_156),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_4),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_73),
.C(n_58),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_146),
.C(n_144),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_162),
.B(n_155),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_143),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_148),
.B(n_12),
.Y(n_163)
);

AOI31xp67_ASAP7_75t_SL g167 ( 
.A1(n_163),
.A2(n_5),
.A3(n_6),
.B(n_9),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.C(n_5),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_160),
.B(n_165),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_10),
.B(n_52),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_166),
.B(n_11),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);


endmodule