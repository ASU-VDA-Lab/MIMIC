module real_jpeg_22530_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_22),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_55),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_2),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_119),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_119),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_119),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_22),
.B1(n_25),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_124),
.Y(n_177)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_131),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_6),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_7),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_9),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_14),
.B(n_47),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_122),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_9),
.A2(n_96),
.B1(n_177),
.B2(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_76),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_29),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_29),
.B(n_206),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_11),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_22),
.B1(n_25),
.B2(n_117),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_117),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_117),
.Y(n_195)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_20),
.A2(n_53),
.B(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_21),
.Y(n_302)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_27),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_22),
.B(n_122),
.CON(n_121),
.SN(n_121)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_31),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_26),
.A2(n_33),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_27),
.B(n_29),
.Y(n_128)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_28),
.A2(n_34),
.B1(n_121),
.B2(n_128),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_28),
.A2(n_41),
.A3(n_66),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_29),
.A2(n_63),
.B(n_64),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_30),
.A2(n_54),
.B(n_58),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_33),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_74),
.C(n_78),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_37),
.A2(n_38),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_51),
.C(n_59),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_39),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_39),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_39),
.A2(n_59),
.B1(n_60),
.B2(n_314),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_45),
.B(n_49),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_40),
.A2(n_49),
.B(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_40),
.A2(n_45),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_40),
.A2(n_45),
.B1(n_173),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_40),
.A2(n_45),
.B1(n_195),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_40),
.A2(n_213),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_40),
.A2(n_45),
.B1(n_104),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_40),
.A2(n_112),
.B(n_248),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_42),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_42),
.A2(n_48),
.B(n_122),
.C(n_169),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_42),
.B(n_64),
.Y(n_207)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_45),
.B(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_46),
.B(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_50),
.B(n_113),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_51),
.A2(n_52),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_58),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_53),
.A2(n_58),
.B1(n_136),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_53),
.A2(n_81),
.B(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_69),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_63),
.A2(n_70),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_63),
.A2(n_70),
.B1(n_116),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_63),
.A2(n_70),
.B1(n_148),
.B2(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_63),
.B(n_73),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_63),
.A2(n_68),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_63),
.A2(n_70),
.B1(n_273),
.B2(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_69),
.A2(n_77),
.B(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_69),
.A2(n_259),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_78),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_331),
.B(n_337),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_307),
.A3(n_326),
.B1(n_329),
.B2(n_330),
.C(n_340),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_286),
.B(n_306),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_264),
.B(n_285),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_153),
.B(n_238),
.C(n_263),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_141),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_90),
.B(n_141),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_125),
.B2(n_140),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_109),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_93),
.B(n_109),
.C(n_140),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_108),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_94),
.B(n_108),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_98),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_102),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_96),
.A2(n_101),
.B1(n_163),
.B2(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_96),
.A2(n_165),
.B(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_96),
.A2(n_97),
.B(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_97),
.B(n_122),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_100),
.A2(n_161),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_105),
.B(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_120),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_126),
.B(n_133),
.C(n_138),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_142),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_147),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_237),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_231),
.B(n_236),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_218),
.B(n_230),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_200),
.B(n_217),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_187),
.B(n_199),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_174),
.B(n_186),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_166),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_170),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_185),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_214),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_220),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_240),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_261),
.B2(n_262),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_249),
.B2(n_250),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_250),
.C(n_262),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_260),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_258),
.C(n_260),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_284),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_277),
.B2(n_278),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_278),
.C(n_284),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_274),
.C(n_276),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_272),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_280),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_297),
.B(n_301),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_282),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_287),
.B(n_288),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_304),
.B2(n_305),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_296),
.C(n_305),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_294),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_309),
.C(n_318),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_295),
.B(n_309),
.CI(n_318),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_301),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_304),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_319),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_319),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_311),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_324),
.C(n_325),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_334),
.Y(n_336)
);


endmodule