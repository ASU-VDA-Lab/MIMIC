module fake_jpeg_4955_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_68)
);

AND2x4_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_18),
.C(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_48),
.B(n_16),
.C(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_34),
.B1(n_23),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_18),
.Y(n_88)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_43),
.B1(n_20),
.B2(n_24),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_62),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_88),
.B1(n_65),
.B2(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_54),
.B1(n_58),
.B2(n_55),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_101),
.B1(n_109),
.B2(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_54),
.B1(n_67),
.B2(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_108),
.B1(n_72),
.B2(n_78),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_55),
.B(n_62),
.C(n_57),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_70),
.B(n_40),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_49),
.B1(n_51),
.B2(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_64),
.C(n_36),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_82),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_16),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_24),
.B(n_70),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_41),
.B1(n_50),
.B2(n_47),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_72),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_109),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_118),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_122),
.B1(n_101),
.B2(n_97),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_85),
.A3(n_24),
.B1(n_78),
.B2(n_63),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_123),
.B(n_129),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_71),
.B1(n_79),
.B2(n_53),
.Y(n_122)
);

OR2x6_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_40),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_43),
.B1(n_87),
.B2(n_83),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_108),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_13),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_50),
.B1(n_41),
.B2(n_27),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_93),
.B1(n_98),
.B2(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_13),
.B(n_1),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_144),
.B(n_154),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_137),
.B1(n_143),
.B2(n_145),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_100),
.B1(n_107),
.B2(n_95),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_123),
.B1(n_14),
.B2(n_2),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_107),
.A3(n_95),
.B1(n_98),
.B2(n_93),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_90),
.B1(n_50),
.B2(n_41),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_90),
.B(n_40),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_153),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_138),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_116),
.B(n_122),
.C(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_26),
.B(n_21),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_158),
.C(n_162),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_123),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_153),
.B(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_118),
.C(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_164),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_126),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_152),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_129),
.C(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_123),
.B1(n_117),
.B2(n_14),
.Y(n_166)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_123),
.B1(n_14),
.B2(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_132),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_0),
.C(n_2),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_0),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_3),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.C(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_3),
.C(n_4),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_187),
.B(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_171),
.B1(n_162),
.B2(n_157),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_197),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_139),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_199),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_150),
.B(n_133),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_161),
.CI(n_170),
.CON(n_204),
.SN(n_204)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_5),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_145),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_4),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_193),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_192),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_215),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_183),
.B(n_193),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_218),
.B(n_8),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_178),
.C(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_219),
.C(n_198),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_191),
.A2(n_160),
.B1(n_157),
.B2(n_7),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_160),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_190),
.B(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_12),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_8),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_180),
.B1(n_181),
.B2(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_5),
.C(n_6),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_223),
.B(n_229),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_202),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_236),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_5),
.C(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_6),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_232),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_219),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_206),
.B1(n_205),
.B2(n_204),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_243),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_246),
.C(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_238),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_8),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_250),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_9),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_9),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_10),
.Y(n_250)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_234),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_221),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_231),
.C(n_235),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_237),
.B(n_238),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_220),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_265),
.B(n_270),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_11),
.B(n_12),
.Y(n_272)
);

NAND2x1p5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_258),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_281),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_254),
.B(n_257),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_263),
.B(n_283),
.C(n_269),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_284),
.B(n_280),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_278),
.B(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_12),
.Y(n_289)
);


endmodule