module fake_jpeg_14565_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_25),
.B1(n_35),
.B2(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_54),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_49),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_4),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_4),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_55),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_7),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_40),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_84),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_103),
.B1(n_27),
.B2(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_38),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_91),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_37),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_104),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_44),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_34),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_21),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_30),
.B(n_29),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_138),
.C(n_142),
.Y(n_145)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_126),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_7),
.B(n_8),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_139),
.B(n_87),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_9),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_132),
.A3(n_76),
.B1(n_98),
.B2(n_15),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_63),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_136),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_29),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_128),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_102),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_63),
.B1(n_32),
.B2(n_11),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_79),
.B1(n_95),
.B2(n_102),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_80),
.B(n_21),
.C(n_10),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_139),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_21),
.B(n_10),
.C(n_11),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_134),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_107),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_82),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_12),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_21),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_12),
.B(n_14),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_66),
.B(n_15),
.C(n_104),
.Y(n_142)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g203 ( 
.A(n_144),
.B(n_149),
.C(n_164),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_152),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_151),
.A2(n_172),
.B1(n_101),
.B2(n_107),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_67),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_73),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_74),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_166),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_92),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_169),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_74),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_70),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_114),
.B(n_70),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_88),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_92),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_88),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_168),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_75),
.B1(n_79),
.B2(n_101),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_123),
.B1(n_136),
.B2(n_75),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_159),
.B1(n_170),
.B2(n_165),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_138),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_192),
.C(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_142),
.C(n_140),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_71),
.C(n_82),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_172),
.B1(n_140),
.B2(n_164),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_118),
.B(n_124),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_190),
.B(n_201),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_149),
.A2(n_125),
.B(n_132),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_112),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_128),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_119),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_151),
.B1(n_156),
.B2(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_137),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_115),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_166),
.B1(n_172),
.B2(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_230)
);

OAI321xp33_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_148),
.A3(n_159),
.B1(n_161),
.B2(n_144),
.C(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_194),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_154),
.B1(n_147),
.B2(n_135),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_183),
.C(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_160),
.B1(n_108),
.B2(n_143),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_223),
.B1(n_186),
.B2(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_108),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_225),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_222),
.B(n_224),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_146),
.B(n_92),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_160),
.B1(n_110),
.B2(n_146),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_72),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_229),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_228),
.C(n_231),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_203),
.C(n_193),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_190),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_236),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_203),
.C(n_193),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_179),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_223),
.B1(n_210),
.B2(n_213),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_177),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_201),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_217),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_207),
.C(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_249),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_208),
.A3(n_220),
.B1(n_215),
.B2(n_207),
.C1(n_222),
.C2(n_206),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_240),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_227),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_209),
.B(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_235),
.B(n_242),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_204),
.B(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_181),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_236),
.B1(n_242),
.B2(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_260),
.B1(n_262),
.B2(n_257),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_261),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_243),
.B1(n_241),
.B2(n_231),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_224),
.B1(n_200),
.B2(n_198),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_267),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_200),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.C(n_268),
.Y(n_271)
);

OAI31xp33_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_218),
.A3(n_202),
.B(n_180),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_263),
.A2(n_262),
.B(n_261),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_260),
.B(n_261),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_267),
.B(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_250),
.C(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_186),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_274),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.Y(n_278)
);


endmodule