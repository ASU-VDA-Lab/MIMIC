module fake_jpeg_21340_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_55),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_17),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_18),
.B(n_34),
.C(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_31),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_29),
.B1(n_34),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_21),
.B1(n_34),
.B2(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_74),
.Y(n_103)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_99),
.B1(n_64),
.B2(n_52),
.Y(n_119)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_18),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_24),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_63),
.CI(n_32),
.CON(n_140),
.SN(n_140)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_45),
.B1(n_36),
.B2(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_27),
.B(n_10),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_112),
.B1(n_62),
.B2(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_54),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_24),
.B(n_28),
.C(n_22),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_86),
.B1(n_97),
.B2(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_103),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_23),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_64),
.C(n_32),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_82),
.C(n_88),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_28),
.B(n_33),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_138),
.B(n_9),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_60),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_79),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_81),
.B(n_99),
.C(n_84),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_85),
.B(n_91),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_60),
.B1(n_59),
.B2(n_71),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_110),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_77),
.A2(n_59),
.B1(n_27),
.B2(n_22),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_101),
.B1(n_107),
.B2(n_111),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_91),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_86),
.B1(n_101),
.B2(n_87),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_158),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_150),
.B(n_153),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_12),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_12),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_115),
.C(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_156),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_85),
.B(n_92),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_131),
.A3(n_122),
.B1(n_138),
.B2(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_161),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_79),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_170),
.B1(n_113),
.B2(n_149),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_23),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_168),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_134),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_11),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_23),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_119),
.C(n_140),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_20),
.B1(n_1),
.B2(n_0),
.Y(n_170)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_176),
.Y(n_215)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_190),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_140),
.B(n_117),
.C(n_135),
.D(n_130),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_192),
.B(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_124),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_170),
.B1(n_161),
.B2(n_149),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_191),
.Y(n_208)
);

NOR4xp25_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_124),
.C(n_127),
.D(n_132),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_132),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_1),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_143),
.B(n_166),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_202),
.B(n_205),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_207),
.C(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_191),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_166),
.B(n_146),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_157),
.B1(n_159),
.B2(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_145),
.B1(n_164),
.B2(n_148),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_155),
.B1(n_167),
.B2(n_142),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_211),
.B1(n_219),
.B2(n_171),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_155),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_150),
.C(n_147),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_160),
.B1(n_151),
.B2(n_139),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_160),
.C(n_20),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_220),
.C(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_3),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_4),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_189),
.B1(n_196),
.B2(n_176),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_3),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_171),
.B1(n_179),
.B2(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_230),
.Y(n_249)
);

XNOR2x2_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_185),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_179),
.B1(n_183),
.B2(n_174),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_186),
.C(n_173),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_205),
.C(n_202),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_186),
.B1(n_182),
.B2(n_7),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_235),
.B1(n_227),
.B2(n_213),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_245),
.C(n_225),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_207),
.C(n_209),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_225),
.C(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_206),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_203),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_210),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_231),
.B(n_228),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_246),
.B1(n_237),
.B2(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_230),
.C(n_234),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_236),
.C(n_199),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_247),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_222),
.C(n_212),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_215),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_269),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_248),
.B1(n_242),
.B2(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.C(n_201),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_254),
.B(n_214),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_277),
.C(n_7),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_268),
.Y(n_279)
);

AOI31xp67_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_216),
.A3(n_255),
.B(n_8),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_4),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_4),
.C(n_7),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_267),
.B(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_281),
.B1(n_8),
.B2(n_11),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_276),
.B(n_11),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_8),
.B(n_14),
.Y(n_286)
);

AOI21x1_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_14),
.B(n_15),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_285),
.C(n_15),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_16),
.B(n_273),
.Y(n_290)
);


endmodule