module fake_jpeg_14819_n_21 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_21);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_21;

wire n_13;
wire n_10;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_0),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_7),
.C(n_9),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_10),
.CI(n_15),
.CON(n_17),
.SN(n_17)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_20),
.A2(n_17),
.B(n_18),
.Y(n_21)
);


endmodule