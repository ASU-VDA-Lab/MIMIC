module fake_jpeg_25872_n_275 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_93;
wire n_54;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_17),
.Y(n_50)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_21),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_41),
.B1(n_43),
.B2(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_61),
.B1(n_62),
.B2(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_64),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_22),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_34),
.B1(n_31),
.B2(n_22),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_40),
.B1(n_36),
.B2(n_44),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_41),
.B(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_32),
.B1(n_19),
.B2(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_68),
.B(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_94),
.B1(n_97),
.B2(n_58),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_39),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_74),
.C(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_77),
.B1(n_95),
.B2(n_100),
.Y(n_103)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_40),
.B1(n_37),
.B2(n_43),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_82),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_40),
.B1(n_36),
.B2(n_63),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_39),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_98),
.C(n_54),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_42),
.B1(n_33),
.B2(n_29),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_66),
.B1(n_46),
.B2(n_56),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_30),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_80),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_56),
.B1(n_24),
.B2(n_54),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_24),
.B1(n_54),
.B2(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_121),
.B1(n_128),
.B2(n_100),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_58),
.B1(n_1),
.B2(n_3),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_134),
.Y(n_170)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_141),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_124),
.B(n_120),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_123),
.B(n_120),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_143),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_147),
.B1(n_158),
.B2(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_70),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_148),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_151),
.C(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_68),
.B1(n_71),
.B2(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_102),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_108),
.B(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_74),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_74),
.C(n_73),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_73),
.C(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_173),
.B1(n_181),
.B2(n_76),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_184),
.B(n_3),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_161),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_168),
.B(n_149),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_105),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_169),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_118),
.B(n_112),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_112),
.B1(n_125),
.B2(n_87),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_88),
.B1(n_94),
.B2(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_89),
.CI(n_98),
.CON(n_176),
.SN(n_176)
);

AOI221xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_156),
.B1(n_146),
.B2(n_130),
.C(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_140),
.B1(n_143),
.B2(n_134),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_98),
.C(n_106),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_154),
.C(n_106),
.Y(n_191)
);

NAND2xp67_ASAP7_75t_SL g184 ( 
.A(n_133),
.B(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_198),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_139),
.C(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_196),
.B(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_200),
.C(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_131),
.B1(n_157),
.B2(n_99),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_195),
.B1(n_206),
.B2(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_6),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_202),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_6),
.C(n_7),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_15),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_167),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_7),
.C(n_8),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_160),
.A3(n_161),
.B1(n_163),
.B2(n_175),
.C1(n_176),
.C2(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_209),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_212),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_169),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_173),
.B(n_177),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_225),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_224),
.B1(n_202),
.B2(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_174),
.B1(n_185),
.B2(n_164),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_174),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_191),
.C(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_230),
.C(n_236),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_192),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_205),
.C(n_200),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_219),
.B1(n_176),
.B2(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_193),
.C(n_199),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_195),
.C(n_194),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_221),
.C(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_216),
.B1(n_215),
.B2(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_242),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_220),
.B1(n_236),
.B2(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_249),
.B1(n_229),
.B2(n_234),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_246),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_219),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_250),
.B1(n_233),
.B2(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_230),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_216),
.B1(n_215),
.B2(n_164),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_226),
.C(n_227),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_258),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_244),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_241),
.B(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_231),
.C(n_196),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_242),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_11),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_268),
.B(n_262),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_258),
.B(n_14),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_268),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_13),
.B(n_14),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.Y(n_275)
);


endmodule