module real_jpeg_7668_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_0),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_0),
.A2(n_22),
.B1(n_65),
.B2(n_68),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_0),
.A2(n_22),
.B1(n_47),
.B2(n_48),
.Y(n_267)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_57),
.B1(n_65),
.B2(n_68),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_4),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_65),
.B1(n_68),
.B2(n_104),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_104),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_104),
.Y(n_222)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_5),
.A2(n_48),
.B(n_60),
.C(n_89),
.D(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_5),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_110),
.B(n_112),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_31),
.B(n_42),
.C(n_146),
.D(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_35),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_28),
.B(n_32),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_127),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_6),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_65),
.B1(n_68),
.B2(n_92),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_92),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_7),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_7),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_130),
.B(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_34),
.B1(n_65),
.B2(n_68),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_14),
.A2(n_55),
.B1(n_65),
.B2(n_68),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_15),
.A2(n_65),
.B1(n_68),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_15),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_109),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_109),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_109),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_16),
.A2(n_65),
.B1(n_68),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_16),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_158),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_158),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_16),
.A2(n_23),
.B1(n_24),
.B2(n_158),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_78),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_25),
.B1(n_35),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_27),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_23),
.A2(n_27),
.B(n_127),
.C(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_25),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_25),
.B(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_26),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_26),
.A2(n_30),
.B1(n_222),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_26),
.A2(n_207),
.B(n_245),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_26),
.A2(n_30),
.B1(n_54),
.B2(n_288),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_30),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_30),
.A2(n_223),
.B(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_35),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_71),
.C(n_73),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_37),
.A2(n_38),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_313),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_50),
.B1(n_167),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_41),
.A2(n_202),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_46),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_42),
.A2(n_46),
.B1(n_242),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_42),
.A2(n_46),
.B1(n_260),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_44),
.B(n_47),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_45),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_48),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_50),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_50),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_50),
.A2(n_168),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_52),
.A2(n_53),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_58),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_69),
.B1(n_103),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_59),
.A2(n_144),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_59),
.A2(n_69),
.B1(n_199),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_59),
.A2(n_69),
.B1(n_217),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_59),
.A2(n_69),
.B1(n_236),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_60),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_60),
.A2(n_64),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_68),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_65),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_111),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_68),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_69),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_69),
.A2(n_105),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_70),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_71),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_331),
.B(n_337),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_304),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_339),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_252),
.A3(n_292),
.B1(n_298),
.B2(n_303),
.C(n_340),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_210),
.C(n_249),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_182),
.B(n_209),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_161),
.B(n_181),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_138),
.B(n_160),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_115),
.B(n_137),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_102),
.C(n_107),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_110),
.A2(n_111),
.B1(n_157),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_110),
.A2(n_111),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_110),
.A2(n_111),
.B1(n_192),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_110),
.A2(n_111),
.B1(n_215),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_110),
.A2(n_111),
.B(n_234),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_119),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_127),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_124),
.B(n_136),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B(n_135),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_128),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_151),
.B2(n_159),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_150),
.C(n_159),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_155),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_178),
.C(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_176),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_195),
.C(n_196),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_191),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_211),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_229),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_229),
.Y(n_301)
);

FAx1_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.CI(n_219),
.CON(n_212),
.SN(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_247),
.B2(n_248),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_237),
.C(n_248),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_243),
.C(n_246),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_251),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_270),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_253),
.B(n_270),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.C(n_269),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_254),
.A2(n_255),
.B1(n_263),
.B2(n_297),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_263),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_265),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_283),
.B(n_287),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_267),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_290),
.B2(n_291),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_281),
.B2(n_282),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_282),
.C(n_291),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_280),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_280),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_280),
.A2(n_306),
.B1(n_315),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_289),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_317),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_317),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_315),
.C(n_316),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_308),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_313),
.C(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_319),
.C(n_323),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_336),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule