module fake_ariane_2733_n_764 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_764);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_764;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_538;
wire n_352;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_458;
wire n_361;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_18),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_9),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_17),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_7),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_91),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_47),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_73),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_55),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_44),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_102),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_8),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_50),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_100),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_4),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_38),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_75),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_57),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_90),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_18),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_51),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_45),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_7),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_145),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_152),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_145),
.B(n_1),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_3),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx11_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_171),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_4),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_5),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_151),
.B(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_196),
.B1(n_163),
.B2(n_167),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_228),
.Y(n_239)
);

OR2x6_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_188),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_150),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_208),
.B1(n_213),
.B2(n_217),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_181),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_184),
.B1(n_191),
.B2(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_194),
.B1(n_182),
.B2(n_180),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_232),
.A2(n_178),
.B1(n_176),
.B2(n_174),
.Y(n_252)
);

CKINVDCx6p67_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_173),
.B1(n_172),
.B2(n_170),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g256 ( 
.A1(n_202),
.A2(n_165),
.B1(n_164),
.B2(n_162),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_160),
.B1(n_157),
.B2(n_10),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_8),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_R g263 ( 
.A1(n_229),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_266)
);

OR2x6_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_12),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_202),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_203),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_271)
);

AO22x2_ASAP7_75t_L g272 ( 
.A1(n_206),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_220),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_214),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_219),
.A2(n_225),
.B1(n_229),
.B2(n_227),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_233),
.A2(n_236),
.B1(n_227),
.B2(n_209),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_231),
.B1(n_221),
.B2(n_218),
.Y(n_280)
);

CKINVDCx6p67_ASAP7_75t_R g281 ( 
.A(n_218),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_236),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_221),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_214),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_260),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_250),
.B(n_236),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_221),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_239),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_224),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_256),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_231),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_240),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_240),
.B(n_224),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_252),
.B(n_235),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

NAND2x1p5_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_218),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_197),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_272),
.B(n_224),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_245),
.B(n_231),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_263),
.B(n_223),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_235),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_241),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_238),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_238),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_223),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_318),
.B(n_235),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_226),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_230),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_285),
.B(n_230),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_226),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_315),
.Y(n_355)
);

OR2x6_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_230),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_226),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_288),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_313),
.A2(n_197),
.B(n_235),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_287),
.B(n_235),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_230),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_226),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_292),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_230),
.Y(n_369)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_197),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_316),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_197),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_324),
.B(n_235),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_292),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_291),
.A2(n_211),
.B(n_210),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_205),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_317),
.B(n_205),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_205),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_293),
.A2(n_211),
.B(n_210),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_298),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_205),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_287),
.B(n_205),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_210),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_284),
.B(n_210),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_299),
.B(n_210),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_314),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_284),
.B(n_330),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g394 ( 
.A(n_290),
.B(n_35),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

OR2x2_ASAP7_75t_SL g396 ( 
.A(n_341),
.B(n_36),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_340),
.B(n_210),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_337),
.B(n_37),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_211),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_294),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_346),
.A2(n_347),
.B(n_290),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_304),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_323),
.B(n_211),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_302),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_329),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_332),
.B(n_211),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_335),
.A2(n_211),
.B(n_41),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_307),
.B(n_40),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_322),
.B(n_142),
.Y(n_415)
);

OR2x6_ASAP7_75t_L g416 ( 
.A(n_414),
.B(n_342),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_342),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_320),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_297),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_331),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_328),
.Y(n_424)
);

NAND2x1_ASAP7_75t_L g425 ( 
.A(n_365),
.B(n_301),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_370),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_359),
.B(n_335),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_372),
.B(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

BUFx4f_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_371),
.B(n_343),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_371),
.B(n_305),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_306),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_356),
.B(n_326),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_309),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

NAND2x1p5_ASAP7_75t_L g444 ( 
.A(n_365),
.B(n_382),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_356),
.B(n_326),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_364),
.B(n_311),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_312),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

NAND2x1p5_ASAP7_75t_L g451 ( 
.A(n_365),
.B(n_308),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_348),
.B(n_310),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_356),
.B(n_310),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_355),
.B(n_42),
.Y(n_454)
);

BUFx8_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_408),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_394),
.B(n_43),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_360),
.B(n_46),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_348),
.B(n_48),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_387),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_358),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_354),
.B(n_381),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_410),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_471),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_394),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_404),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_460),
.A2(n_398),
.B1(n_399),
.B2(n_402),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_429),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_398),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_419),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_419),
.Y(n_488)
);

CKINVDCx6p67_ASAP7_75t_R g489 ( 
.A(n_416),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_424),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_433),
.B(n_399),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_455),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_433),
.B(n_381),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_433),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_416),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_385),
.Y(n_502)
);

BUFx5_ASAP7_75t_L g503 ( 
.A(n_430),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_456),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_456),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_416),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_514),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_509),
.Y(n_520)
);

BUFx8_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_420),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

BUFx6f_ASAP7_75t_SL g525 ( 
.A(n_491),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_485),
.A2(n_422),
.B1(n_420),
.B2(n_445),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_479),
.A2(n_466),
.B(n_473),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_479),
.A2(n_396),
.B1(n_442),
.B2(n_434),
.Y(n_528)
);

BUFx2_ASAP7_75t_SL g529 ( 
.A(n_491),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_476),
.A2(n_396),
.B1(n_457),
.B2(n_432),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_480),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_480),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_476),
.A2(n_461),
.B1(n_492),
.B2(n_498),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_483),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_478),
.A2(n_440),
.B1(n_445),
.B2(n_422),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_517),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_483),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_494),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_501),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_492),
.A2(n_459),
.B1(n_467),
.B2(n_472),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_503),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_474),
.A2(n_440),
.B1(n_445),
.B2(n_412),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_492),
.A2(n_420),
.B1(n_423),
.B2(n_401),
.Y(n_546)
);

AOI21xp33_ASAP7_75t_L g547 ( 
.A1(n_478),
.A2(n_363),
.B(n_437),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_492),
.A2(n_423),
.B1(n_401),
.B2(n_448),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_493),
.A2(n_415),
.B1(n_439),
.B2(n_413),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_502),
.B(n_459),
.Y(n_550)
);

CKINVDCx11_ASAP7_75t_R g551 ( 
.A(n_490),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_513),
.A2(n_472),
.B1(n_467),
.B2(n_438),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_481),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

INVx6_ASAP7_75t_SL g555 ( 
.A(n_489),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_502),
.A2(n_423),
.B1(n_439),
.B2(n_469),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_500),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_491),
.Y(n_559)
);

BUFx2_ASAP7_75t_SL g560 ( 
.A(n_505),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_520),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_SL g562 ( 
.A1(n_530),
.A2(n_528),
.B1(n_549),
.B2(n_534),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_530),
.B(n_503),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_528),
.A2(n_505),
.B1(n_499),
.B2(n_503),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_550),
.A2(n_454),
.B1(n_402),
.B2(n_499),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_511),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_534),
.A2(n_505),
.B1(n_511),
.B2(n_518),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g570 ( 
.A1(n_527),
.A2(n_369),
.B(n_362),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_386),
.B(n_373),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_554),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_544),
.A2(n_386),
.B1(n_511),
.B2(n_489),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_526),
.A2(n_402),
.B1(n_501),
.B2(n_508),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_523),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_532),
.B(n_501),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_501),
.B1(n_508),
.B2(n_382),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_552),
.A2(n_503),
.B1(n_518),
.B2(n_515),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_536),
.A2(n_551),
.B1(n_542),
.B2(n_546),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_559),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_542),
.A2(n_503),
.B1(n_518),
.B2(n_515),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_536),
.A2(n_518),
.B1(n_439),
.B2(n_484),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_547),
.A2(n_518),
.B1(n_497),
.B2(n_507),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_524),
.B(n_518),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_519),
.B(n_521),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_521),
.B(n_503),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_547),
.A2(n_495),
.B1(n_512),
.B2(n_484),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_537),
.A2(n_501),
.B1(n_508),
.B2(n_464),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_525),
.A2(n_557),
.B1(n_545),
.B2(n_560),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_533),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_556),
.B(n_380),
.C(n_385),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_558),
.A2(n_508),
.B(n_486),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_543),
.A2(n_508),
.B1(n_496),
.B2(n_510),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_503),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_541),
.A2(n_507),
.B1(n_495),
.B2(n_512),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_529),
.A2(n_486),
.B1(n_510),
.B2(n_496),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_538),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_380),
.C(n_452),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_525),
.A2(n_515),
.B1(n_503),
.B2(n_446),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_553),
.A2(n_497),
.B1(n_515),
.B2(n_516),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_545),
.A2(n_496),
.B1(n_486),
.B2(n_510),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_557),
.B(n_477),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_558),
.A2(n_503),
.B1(n_515),
.B2(n_447),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_591),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_562),
.A2(n_565),
.B1(n_579),
.B2(n_581),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_562),
.A2(n_465),
.B1(n_468),
.B2(n_462),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_565),
.A2(n_486),
.B1(n_496),
.B2(n_510),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_494),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_SL g613 ( 
.A(n_601),
.B(n_540),
.C(n_389),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_592),
.A2(n_516),
.B1(n_506),
.B2(n_462),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_571),
.A2(n_465),
.B1(n_468),
.B2(n_405),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_567),
.A2(n_506),
.B1(n_540),
.B2(n_488),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_581),
.A2(n_487),
.B1(n_555),
.B2(n_458),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_574),
.A2(n_487),
.B1(n_488),
.B2(n_482),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_482),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_590),
.B(n_599),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_578),
.A2(n_555),
.B1(n_458),
.B2(n_427),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_577),
.A2(n_488),
.B1(n_482),
.B2(n_361),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_569),
.A2(n_441),
.B1(n_397),
.B2(n_391),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_578),
.A2(n_397),
.B1(n_395),
.B2(n_391),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_576),
.A2(n_358),
.B1(n_389),
.B2(n_352),
.Y(n_625)
);

AO22x1_ASAP7_75t_L g626 ( 
.A1(n_580),
.A2(n_458),
.B1(n_427),
.B2(n_351),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_564),
.A2(n_427),
.B1(n_444),
.B2(n_367),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_586),
.A2(n_444),
.B1(n_367),
.B2(n_426),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_582),
.A2(n_397),
.B1(n_395),
.B2(n_391),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_573),
.A2(n_391),
.B1(n_395),
.B2(n_406),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_593),
.B(n_367),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_583),
.A2(n_391),
.B1(n_395),
.B2(n_406),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_563),
.A2(n_395),
.B1(n_406),
.B2(n_407),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_589),
.A2(n_426),
.B1(n_388),
.B2(n_411),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_566),
.A2(n_587),
.B1(n_588),
.B2(n_603),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_602),
.A2(n_388),
.B1(n_411),
.B2(n_349),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_607),
.A2(n_451),
.B1(n_384),
.B2(n_425),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_561),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_570),
.A2(n_406),
.B1(n_374),
.B2(n_384),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_606),
.B(n_366),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_580),
.A2(n_406),
.B1(n_390),
.B2(n_451),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_607),
.B(n_378),
.C(n_377),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_608),
.B(n_585),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_572),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_596),
.Y(n_645)
);

AOI211xp5_ASAP7_75t_L g646 ( 
.A1(n_609),
.A2(n_605),
.B(n_594),
.C(n_604),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_626),
.B(n_572),
.C(n_561),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_612),
.B(n_584),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_619),
.B(n_595),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_610),
.A2(n_598),
.B(n_597),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_638),
.B(n_366),
.Y(n_651)
);

OAI21xp33_ASAP7_75t_L g652 ( 
.A1(n_610),
.A2(n_377),
.B(n_366),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_640),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_616),
.B(n_377),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_639),
.C(n_631),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_617),
.B(n_377),
.Y(n_656)
);

AOI221xp5_ASAP7_75t_L g657 ( 
.A1(n_615),
.A2(n_383),
.B1(n_376),
.B2(n_377),
.C(n_56),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_615),
.B(n_621),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_618),
.B(n_141),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_624),
.B(n_49),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_625),
.A2(n_52),
.B(n_54),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_611),
.B(n_139),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_58),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_138),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_641),
.B(n_59),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_SL g666 ( 
.A1(n_634),
.A2(n_614),
.B1(n_642),
.B2(n_623),
.C(n_630),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_627),
.B(n_60),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_622),
.B(n_62),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_63),
.Y(n_669)
);

AOI221xp5_ASAP7_75t_L g670 ( 
.A1(n_633),
.A2(n_629),
.B1(n_636),
.B2(n_632),
.C(n_67),
.Y(n_670)
);

OR2x6_ASAP7_75t_SL g671 ( 
.A(n_655),
.B(n_64),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_65),
.Y(n_672)
);

NAND2x1_ASAP7_75t_L g673 ( 
.A(n_643),
.B(n_66),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_648),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_645),
.B(n_68),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_661),
.B(n_69),
.C(n_70),
.Y(n_677)
);

OR2x2_ASAP7_75t_SL g678 ( 
.A(n_658),
.B(n_649),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_670),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_651),
.B(n_78),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_650),
.B(n_654),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_656),
.Y(n_683)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_644),
.B(n_79),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_669),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_651),
.B(n_85),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_678),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_681),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_683),
.B(n_647),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_675),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_682),
.B(n_646),
.Y(n_691)
);

XOR2x2_ASAP7_75t_L g692 ( 
.A(n_677),
.B(n_666),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_674),
.B(n_686),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_676),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_669),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_672),
.Y(n_696)
);

AND4x1_ASAP7_75t_L g697 ( 
.A(n_677),
.B(n_668),
.C(n_662),
.D(n_665),
.Y(n_697)
);

XOR2x2_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_684),
.Y(n_698)
);

NOR2x1_ASAP7_75t_R g699 ( 
.A(n_691),
.B(n_671),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_688),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_694),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_690),
.Y(n_702)
);

OAI22x1_ASAP7_75t_L g703 ( 
.A1(n_702),
.A2(n_687),
.B1(n_691),
.B2(n_697),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_701),
.A2(n_689),
.B1(n_696),
.B2(n_695),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_700),
.Y(n_705)
);

OA22x2_ASAP7_75t_L g706 ( 
.A1(n_698),
.A2(n_695),
.B1(n_689),
.B2(n_692),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_705),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_703),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_709),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_709),
.A2(n_706),
.B1(n_699),
.B2(n_700),
.Y(n_711)
);

NAND4xp75_ASAP7_75t_L g712 ( 
.A(n_708),
.B(n_685),
.C(n_676),
.D(n_663),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_710),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_712),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_SL g715 ( 
.A1(n_711),
.A2(n_707),
.B(n_673),
.C(n_697),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_710),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_713),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_716),
.A2(n_696),
.B1(n_693),
.B2(n_665),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_714),
.A2(n_679),
.B1(n_693),
.B2(n_660),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_715),
.B(n_659),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_715),
.Y(n_721)
);

NOR4xp25_ASAP7_75t_L g722 ( 
.A(n_716),
.B(n_679),
.C(n_664),
.D(n_667),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_716),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_717),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_722),
.B(n_667),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_719),
.A2(n_660),
.B1(n_652),
.B2(n_657),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_718),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_720),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_725),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_729),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_727),
.Y(n_733)
);

AND5x1_ASAP7_75t_L g734 ( 
.A(n_724),
.B(n_86),
.C(n_87),
.D(n_88),
.E(n_89),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_726),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_728),
.Y(n_737)
);

AND4x1_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_97),
.C(n_98),
.D(n_99),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_725),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_739),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_731),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_732),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_736),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_733),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_737),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_734),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_742),
.A2(n_738),
.B1(n_103),
.B2(n_104),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_101),
.B1(n_105),
.B2(n_107),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_746),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_750)
);

OAI22x1_ASAP7_75t_L g751 ( 
.A1(n_740),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_741),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_752),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_750),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_743),
.B1(n_744),
.B2(n_745),
.Y(n_757)
);

NAND4xp25_ASAP7_75t_L g758 ( 
.A(n_755),
.B(n_743),
.C(n_749),
.D(n_121),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_118),
.B1(n_120),
.B2(n_123),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_757),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_758),
.B1(n_759),
.B2(n_756),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_761),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_762),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.C(n_129),
.Y(n_763)
);

AOI211xp5_ASAP7_75t_L g764 ( 
.A1(n_763),
.A2(n_131),
.B(n_134),
.C(n_135),
.Y(n_764)
);


endmodule