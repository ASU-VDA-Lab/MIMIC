module real_jpeg_17981_n_23 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_51;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_62),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_1),
.B(n_54),
.C(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_2),
.A2(n_25),
.B1(n_57),
.B2(n_58),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_57),
.B1(n_64),
.B2(n_83),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_17),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.C(n_82),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_4),
.B(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_6),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_38),
.C(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.C(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_21),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_72),
.C(n_81),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_14),
.B(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_44),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_47),
.C(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp67_ASAP7_75t_SL g66 ( 
.A(n_16),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_18),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

AOI222xp33_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_24),
.B1(n_59),
.B2(n_63),
.C1(n_84),
.C2(n_86),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B(n_56),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_52),
.B(n_55),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_50),
.B(n_51),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_46),
.B(n_49),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_44),
.C(n_45),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B(n_43),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_42),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B(n_80),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);


endmodule