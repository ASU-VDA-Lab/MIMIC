module fake_jpeg_144_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_18),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_35),
.B(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_1),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_20),
.B1(n_22),
.B2(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_67),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_20),
.B1(n_17),
.B2(n_21),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_66),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_34),
.A2(n_29),
.B1(n_19),
.B2(n_18),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_29),
.C(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_1),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_51),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_36),
.A2(n_32),
.B1(n_16),
.B2(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_44),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_49),
.B1(n_44),
.B2(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_76),
.B1(n_54),
.B2(n_68),
.Y(n_108)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_37),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_73),
.B(n_7),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_103),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_5),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_53),
.B1(n_55),
.B2(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_73),
.B1(n_58),
.B2(n_79),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_73),
.B1(n_79),
.B2(n_6),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_102),
.B(n_92),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_100),
.B1(n_93),
.B2(n_90),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_6),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_84),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.C(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_88),
.C(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_115),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_98),
.C(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_116),
.B1(n_122),
.B2(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_113),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_87),
.B(n_79),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_137),
.A2(n_127),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_141),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_119),
.C(n_117),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_115),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_134),
.C(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_158),
.B(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_124),
.B1(n_123),
.B2(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_154),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_117),
.A3(n_136),
.B1(n_118),
.B2(n_121),
.C1(n_126),
.C2(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_144),
.C(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_129),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_142),
.B(n_148),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_157),
.B(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_164),
.C(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_144),
.C(n_146),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_152),
.A3(n_153),
.B1(n_139),
.B2(n_156),
.C1(n_136),
.C2(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_159),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_162),
.C(n_106),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_173),
.B(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_114),
.B(n_107),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_79),
.Y(n_177)
);


endmodule