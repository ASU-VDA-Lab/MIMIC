module real_jpeg_7918_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_320, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_320;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_1),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_36),
.B1(n_49),
.B2(n_52),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_4),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_143),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_49),
.B1(n_52),
.B2(n_143),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_143),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_10),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_49),
.B1(n_52),
.B2(n_161),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_161),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_161),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_49),
.B1(n_52),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_13),
.A2(n_49),
.B1(n_52),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_170),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_170),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_170),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_14),
.A2(n_33),
.B1(n_49),
.B2(n_52),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_14),
.A2(n_33),
.B1(n_66),
.B2(n_67),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_15),
.A2(n_52),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_15),
.B(n_52),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_15),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_15),
.A2(n_90),
.B1(n_93),
.B2(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_15),
.B(n_105),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_15),
.A2(n_25),
.B(n_27),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_179),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_86),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_21),
.A2(n_74),
.B1(n_75),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_21),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_22),
.A2(n_23),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_60),
.C(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_29),
.B(n_32),
.C(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_24),
.A2(n_38),
.B1(n_262),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_24),
.A2(n_38),
.B1(n_142),
.B2(n_271),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_45),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g204 ( 
.A(n_27),
.B(n_179),
.CON(n_204),
.SN(n_204)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_29),
.A2(n_32),
.B(n_179),
.C(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_35),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_37),
.A2(n_105),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_38),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_38),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_53),
.B(n_56),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_43),
.A2(n_59),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_43),
.A2(n_59),
.B1(n_222),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_43),
.A2(n_115),
.B(n_258),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_48),
.B1(n_54),
.B2(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_44),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_44),
.A2(n_48),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_44),
.A2(n_57),
.B(n_116),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_45),
.B(n_52),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_49),
.B1(n_204),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_48),
.B(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_78),
.B(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_59),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_61),
.B1(n_114),
.B2(n_119),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_70),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_65),
.B1(n_97),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_65),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_62),
.A2(n_65),
.B1(n_169),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_62),
.A2(n_65),
.B1(n_194),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_62),
.A2(n_80),
.B(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_65),
.B(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_65),
.A2(n_82),
.B(n_139),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_66),
.B(n_69),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_66),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_67),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_71),
.A2(n_85),
.B(n_99),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_86),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_100),
.B(n_101),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_100),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_89),
.A2(n_96),
.B1(n_100),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_90),
.A2(n_93),
.B1(n_160),
.B2(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_90),
.A2(n_137),
.B(n_163),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_90),
.A2(n_94),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_90),
.A2(n_93),
.B1(n_226),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_90),
.A2(n_212),
.B(n_248),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_91),
.A2(n_92),
.B1(n_159),
.B2(n_162),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_92),
.B(n_136),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_179),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_93),
.A2(n_135),
.B(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_96),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_121),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_120),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_150),
.B(n_318),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_147),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_125),
.B(n_147),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_126),
.B(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_126),
.B(n_310),
.Y(n_317)
);

FAx1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.CI(n_132),
.CON(n_126),
.SN(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.C(n_145),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_133),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_134),
.B(n_138),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_297),
.A3(n_309),
.B1(n_311),
.B2(n_317),
.C(n_320),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_264),
.C(n_293),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_238),
.B(n_263),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_215),
.B(n_237),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_197),
.B(n_214),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_188),
.B(n_196),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_176),
.B(n_187),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_171),
.B2(n_175),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_175),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_171),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_182),
.B(n_186),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_198),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_193),
.CI(n_195),
.CON(n_191),
.SN(n_191)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_208),
.B2(n_213),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_207),
.C(n_213),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_231),
.B2(n_232),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_234),
.C(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_230),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_240),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_252),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_251),
.C(n_252),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_280),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_280),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_274),
.C(n_278),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_269),
.C(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_289),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_285),
.C(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_312),
.B(n_316),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_300),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_306),
.C(n_308),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B(n_315),
.Y(n_312)
);


endmodule