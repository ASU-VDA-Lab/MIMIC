module fake_netlist_6_2078_n_1435 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1435);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1435;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx2_ASAP7_75t_L g329 ( 
.A(n_110),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_289),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_179),
.B(n_303),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_124),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_210),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_82),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_61),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_234),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_128),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_72),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_25),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_145),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_235),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_240),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_172),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_10),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_135),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_43),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_286),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_14),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_22),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_299),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_58),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_174),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_79),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_308),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_23),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_0),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_224),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_305),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_229),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_87),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_215),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_134),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_33),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_232),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_68),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_249),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_157),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_38),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_143),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_21),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_270),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_221),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_85),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_129),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_194),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_13),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_96),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_141),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_130),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_20),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_244),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_120),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_230),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_245),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_25),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_231),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_24),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_105),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_152),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_204),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_119),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_165),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_39),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_40),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_153),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_181),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_15),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_131),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_288),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_239),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_252),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_164),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_212),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_171),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_24),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_81),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_35),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_142),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_185),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_320),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_63),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_326),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_139),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_104),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_14),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_90),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_168),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_74),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_156),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_149),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_19),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_187),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_297),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_191),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_264),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_2),
.Y(n_443)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_247),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_121),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_140),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_290),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_114),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_76),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_66),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_163),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_293),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_176),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_274),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_127),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_267),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_89),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_315),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_88),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_51),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_195),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_31),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_225),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_217),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_57),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_55),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_77),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_159),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_298),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_222),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_32),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_23),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_256),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_192),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_107),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_102),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_220),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_287),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_155),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_100),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_59),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_126),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_189),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_322),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_246),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_43),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_0),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_227),
.Y(n_488)
);

HB1xp67_ASAP7_75t_SL g489 ( 
.A(n_92),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_291),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_312),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_273),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_50),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_93),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_266),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_84),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_98),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_251),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_248),
.B(n_86),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_42),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_117),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_170),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_276),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_37),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_151),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_147),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_216),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_238),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_205),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_213),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_219),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_28),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_292),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_199),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_83),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_133),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_259),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_28),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_254),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_111),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_209),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_203),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_45),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_226),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_73),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_309),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_175),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_241),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_173),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_132),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_67),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_328),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_33),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_233),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_53),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_103),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_243),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_21),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_323),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_8),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_186),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_284),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_311),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_190),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_177),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_65),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_64),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_381),
.Y(n_548)
);

AOI22x1_ASAP7_75t_SL g549 ( 
.A1(n_379),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_365),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

BUFx12f_ASAP7_75t_L g554 ( 
.A(n_381),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_357),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_373),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_398),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_3),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_366),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_330),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_385),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_385),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_373),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_478),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_518),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_385),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_385),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_348),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_444),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_459),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_459),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_400),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_351),
.B(n_4),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_355),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_467),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_4),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_358),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_418),
.B(n_5),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_374),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_332),
.A2(n_335),
.B(n_334),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_546),
.B(n_5),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_467),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_352),
.B(n_6),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_387),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_484),
.B(n_7),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_391),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_486),
.Y(n_595)
);

OA21x2_ASAP7_75t_L g596 ( 
.A1(n_337),
.A2(n_9),
.B(n_11),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_347),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_410),
.Y(n_598)
);

CKINVDCx6p67_ASAP7_75t_R g599 ( 
.A(n_364),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_484),
.B(n_46),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_437),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_333),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

AOI22x1_ASAP7_75t_SL g604 ( 
.A1(n_407),
.A2(n_443),
.B1(n_471),
.B2(n_462),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_333),
.B(n_12),
.Y(n_605)
);

AOI22x1_ASAP7_75t_SL g606 ( 
.A1(n_487),
.A2(n_500),
.B1(n_512),
.B2(n_504),
.Y(n_606)
);

BUFx8_ASAP7_75t_L g607 ( 
.A(n_353),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_533),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_362),
.B(n_12),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_467),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_329),
.A2(n_48),
.B(n_47),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_390),
.B(n_15),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_362),
.B(n_16),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_456),
.B(n_16),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_444),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_342),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_392),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_488),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_370),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_537),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_540),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_382),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_537),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_456),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_393),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_453),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_336),
.B(n_17),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_532),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_340),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_375),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_345),
.Y(n_635)
);

INVx6_ASAP7_75t_L g636 ( 
.A(n_479),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_346),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_376),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_430),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_479),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_338),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_523),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_479),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_479),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_413),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_409),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_349),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_434),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g649 ( 
.A(n_339),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_419),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_419),
.B(n_27),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_354),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_352),
.B(n_361),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_454),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_457),
.A2(n_52),
.B(n_49),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_341),
.Y(n_657)
);

OAI22x1_ASAP7_75t_SL g658 ( 
.A1(n_404),
.A2(n_415),
.B1(n_435),
.B2(n_432),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_524),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_371),
.B(n_29),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_372),
.A2(n_56),
.B(n_54),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_380),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_389),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_394),
.Y(n_664)
);

BUFx8_ASAP7_75t_SL g665 ( 
.A(n_438),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_396),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_479),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_397),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_411),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_343),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_403),
.B(n_29),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_344),
.Y(n_672)
);

CKINVDCx6p67_ASAP7_75t_R g673 ( 
.A(n_450),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_416),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_417),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_506),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_427),
.Y(n_677)
);

NOR2x1_ASAP7_75t_L g678 ( 
.A(n_499),
.B(n_60),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_489),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_440),
.B(n_30),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_446),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

OAI22x1_ASAP7_75t_L g683 ( 
.A1(n_447),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_683)
);

BUFx12f_ASAP7_75t_L g684 ( 
.A(n_350),
.Y(n_684)
);

BUFx8_ASAP7_75t_L g685 ( 
.A(n_331),
.Y(n_685)
);

INVx6_ASAP7_75t_L g686 ( 
.A(n_356),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_451),
.B(n_34),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_455),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_359),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_360),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_448),
.B(n_34),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_458),
.B(n_35),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_461),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_476),
.B(n_36),
.Y(n_694)
);

AND3x2_ASAP7_75t_L g695 ( 
.A(n_578),
.B(n_692),
.C(n_691),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_R g696 ( 
.A(n_571),
.B(n_36),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_665),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_561),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_672),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_602),
.B(n_545),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_553),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_562),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_553),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_619),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_562),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_563),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_690),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_622),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_679),
.B(n_463),
.Y(n_712)
);

CKINVDCx16_ASAP7_75t_R g713 ( 
.A(n_676),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_684),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_673),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_599),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_670),
.B(n_363),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_685),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_641),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_620),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_657),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_575),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_639),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_598),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_624),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_620),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_686),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_679),
.B(n_367),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_576),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_686),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_689),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_580),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_645),
.B(n_474),
.Y(n_734)
);

NOR2xp67_ASAP7_75t_L g735 ( 
.A(n_679),
.B(n_475),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_580),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_590),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_632),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_590),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_689),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_556),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_689),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_548),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_554),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_603),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_603),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_645),
.B(n_481),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_632),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_610),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_R g750 ( 
.A(n_564),
.B(n_368),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_682),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_610),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_658),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_571),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_612),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_612),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_614),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_582),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_608),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_608),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_565),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_642),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_594),
.A2(n_495),
.B1(n_491),
.B2(n_492),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_R g764 ( 
.A(n_596),
.B(n_369),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_570),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_607),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_604),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_623),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_623),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_560),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_574),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_597),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_577),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_625),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_601),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_618),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_551),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_626),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_560),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_606),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_604),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_634),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_654),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_628),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_629),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_630),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_763),
.B(n_581),
.C(n_558),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_700),
.B(n_613),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_762),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_762),
.B(n_585),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_774),
.B(n_671),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_723),
.B(n_630),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_710),
.Y(n_794)
);

BUFx5_ASAP7_75t_L g795 ( 
.A(n_705),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_772),
.B(n_569),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_779),
.B(n_569),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_785),
.B(n_589),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_SL g799 ( 
.A(n_784),
.B(n_621),
.C(n_652),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_704),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_783),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_779),
.B(n_569),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_756),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_774),
.B(n_593),
.C(n_591),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_773),
.B(n_694),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_729),
.B(n_573),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_786),
.B(n_627),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_731),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_733),
.B(n_573),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_737),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_745),
.B(n_573),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_775),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_754),
.B(n_666),
.C(n_663),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_698),
.B(n_631),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_749),
.B(n_755),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_770),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_756),
.B(n_627),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_787),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_756),
.B(n_600),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_756),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_702),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_732),
.B(n_600),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_769),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_740),
.B(n_588),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_758),
.B(n_652),
.C(n_677),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_707),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_717),
.B(n_678),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_708),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_742),
.B(n_588),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_722),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_734),
.B(n_660),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_736),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_706),
.B(n_596),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_739),
.Y(n_834)
);

AOI221xp5_ASAP7_75t_L g835 ( 
.A1(n_759),
.A2(n_683),
.B1(n_680),
.B2(n_595),
.C(n_650),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_760),
.B(n_677),
.C(n_609),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_746),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_747),
.B(n_752),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_720),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_741),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_720),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_695),
.B(n_615),
.C(n_605),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_757),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_766),
.B(n_687),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_701),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_703),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_721),
.B(n_635),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_699),
.B(n_616),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_709),
.B(n_647),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_771),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_712),
.B(n_668),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_735),
.B(n_675),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_761),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_696),
.B(n_552),
.C(n_669),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_711),
.B(n_664),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_728),
.B(n_634),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_750),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_696),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_727),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_765),
.B(n_377),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_716),
.B(n_378),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_730),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_715),
.B(n_633),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_706),
.B(n_383),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_767),
.B(n_384),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_743),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_751),
.B(n_638),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_719),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_697),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_714),
.B(n_638),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_794),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_858),
.B(n_724),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_814),
.B(n_646),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_790),
.B(n_725),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_840),
.B(n_744),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_815),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_792),
.B(n_646),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_808),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_805),
.B(n_386),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_810),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_SL g883 ( 
.A(n_799),
.B(n_782),
.C(n_781),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_843),
.A2(n_494),
.B1(n_496),
.B2(n_490),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_831),
.B(n_648),
.Y(n_885)
);

INVx5_ASAP7_75t_L g886 ( 
.A(n_860),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_800),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_850),
.B(n_388),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_816),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_SL g890 ( 
.A1(n_804),
.A2(n_549),
.B1(n_777),
.B2(n_776),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_824),
.B(n_655),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_829),
.B(n_655),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_826),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_828),
.B(n_579),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_848),
.B(n_659),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_834),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_842),
.B(n_713),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_803),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_795),
.B(n_788),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_846),
.B(n_584),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_793),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_864),
.B(n_395),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_859),
.A2(n_633),
.B(n_653),
.C(n_637),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_860),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_855),
.B(n_835),
.C(n_825),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_860),
.B(n_586),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_801),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_833),
.A2(n_511),
.B1(n_514),
.B2(n_509),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_870),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_854),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_823),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_818),
.B(n_868),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_830),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_847),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_851),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_795),
.B(n_659),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_795),
.B(n_517),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_778),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_849),
.B(n_525),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_854),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_832),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_822),
.A2(n_530),
.B1(n_534),
.B2(n_526),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_856),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_841),
.B(n_726),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_838),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_845),
.A2(n_661),
.B(n_568),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_863),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_827),
.A2(n_789),
.B1(n_791),
.B2(n_836),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_840),
.B(n_867),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_812),
.B(n_399),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_839),
.B(n_796),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_844),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_797),
.B(n_541),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_817),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_802),
.B(n_542),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_803),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_857),
.B(n_543),
.Y(n_938)
);

INVxp33_ASAP7_75t_SL g939 ( 
.A(n_862),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_840),
.B(n_401),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_803),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_837),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_837),
.B(n_555),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_820),
.B(n_637),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_813),
.B(n_402),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_871),
.B(n_405),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_798),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_820),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_861),
.B(n_738),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_820),
.B(n_653),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_865),
.A2(n_412),
.B1(n_414),
.B2(n_408),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_869),
.B(n_592),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_806),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_866),
.A2(n_764),
.B1(n_422),
.B2(n_423),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_807),
.B(n_555),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_809),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_811),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_852),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_853),
.B(n_550),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_932),
.B(n_420),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_891),
.A2(n_656),
.B(n_611),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_892),
.A2(n_583),
.B(n_572),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_926),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_878),
.B(n_424),
.Y(n_964)
);

NOR2x1_ASAP7_75t_L g965 ( 
.A(n_905),
.B(n_748),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_874),
.A2(n_617),
.B(n_587),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_926),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_944),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_919),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_886),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_886),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_900),
.A2(n_426),
.B1(n_428),
.B2(n_425),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_875),
.B(n_429),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_874),
.B(n_431),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_872),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_886),
.B(n_433),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_890),
.A2(n_768),
.B1(n_753),
.B2(n_718),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_880),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_906),
.A2(n_693),
.B(n_662),
.C(n_643),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_939),
.B(n_436),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_902),
.B(n_557),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_921),
.B(n_439),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_882),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_899),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_929),
.A2(n_515),
.B1(n_442),
.B2(n_445),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_904),
.A2(n_693),
.B(n_662),
.C(n_640),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_879),
.B(n_441),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_905),
.B(n_549),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_921),
.B(n_449),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_911),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_958),
.B(n_452),
.Y(n_991)
);

AO32x2_ASAP7_75t_L g992 ( 
.A1(n_923),
.A2(n_37),
.A3(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_887),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_907),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_924),
.B(n_460),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_952),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_899),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_888),
.B(n_464),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_907),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_885),
.A2(n_651),
.B(n_644),
.Y(n_1000)
);

AOI22x1_ASAP7_75t_L g1001 ( 
.A1(n_927),
.A2(n_519),
.B1(n_466),
.B2(n_468),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_935),
.A2(n_520),
.B1(n_469),
.B2(n_470),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_958),
.B(n_465),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_917),
.A2(n_667),
.B(n_477),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_898),
.Y(n_1005)
);

OA21x2_ASAP7_75t_L g1006 ( 
.A1(n_918),
.A2(n_559),
.B(n_557),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_956),
.A2(n_480),
.B(n_473),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_SL g1008 ( 
.A1(n_881),
.A2(n_566),
.B(n_636),
.C(n_674),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_956),
.A2(n_483),
.B(n_482),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_937),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_953),
.A2(n_493),
.B(n_485),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_889),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_957),
.A2(n_498),
.B(n_497),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_922),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_933),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_942),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_920),
.B(n_895),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_950),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_947),
.A2(n_529),
.B1(n_502),
.B2(n_503),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_913),
.B(n_566),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_896),
.B(n_501),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_925),
.B(n_505),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_928),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_938),
.B(n_507),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_909),
.B(n_508),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_899),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_914),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_934),
.A2(n_516),
.B(n_510),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_936),
.A2(n_522),
.B(n_521),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_943),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_910),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_954),
.A2(n_539),
.B1(n_527),
.B2(n_531),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_959),
.A2(n_636),
.B1(n_681),
.B2(n_674),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_941),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_893),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_930),
.B(n_535),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_969),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_963),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_967),
.B(n_912),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1023),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_984),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_961),
.A2(n_916),
.B(n_908),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1006),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_1008),
.A2(n_894),
.B(n_897),
.Y(n_1045)
);

INVx6_ASAP7_75t_SL g1046 ( 
.A(n_990),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_962),
.A2(n_894),
.B(n_915),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_966),
.A2(n_884),
.B(n_903),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_1031),
.Y(n_1049)
);

CKINVDCx8_ASAP7_75t_R g1050 ( 
.A(n_1005),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_984),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_984),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_993),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_999),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1017),
.A2(n_931),
.B(n_946),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_SL g1056 ( 
.A1(n_970),
.A2(n_951),
.B(n_959),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_1016),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_994),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1026),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_987),
.A2(n_945),
.B(n_940),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_1026),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_996),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_997),
.B(n_901),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_960),
.A2(n_959),
.B(n_901),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1001),
.A2(n_873),
.B(n_876),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1014),
.B(n_883),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_1026),
.Y(n_1067)
);

AOI22x1_ASAP7_75t_L g1068 ( 
.A1(n_968),
.A2(n_1018),
.B1(n_1015),
.B2(n_1000),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_1030),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_997),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_971),
.Y(n_1071)
);

INVx6_ASAP7_75t_SL g1072 ( 
.A(n_965),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1034),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_973),
.A2(n_959),
.B(n_955),
.Y(n_1074)
);

AO21x2_ASAP7_75t_L g1075 ( 
.A1(n_991),
.A2(n_955),
.B(n_877),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_1034),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_981),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1027),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1035),
.B(n_62),
.Y(n_1079)
);

INVx3_ASAP7_75t_SL g1080 ( 
.A(n_980),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1006),
.Y(n_1081)
);

INVx3_ASAP7_75t_SL g1082 ( 
.A(n_982),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1034),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_975),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_1003),
.A2(n_949),
.B(n_547),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_983),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_1010),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1012),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1037),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1022),
.B(n_681),
.Y(n_1091)
);

AOI22x1_ASAP7_75t_L g1092 ( 
.A1(n_1020),
.A2(n_544),
.B1(n_536),
.B2(n_688),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1037),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1004),
.A2(n_206),
.B(n_324),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_974),
.A2(n_202),
.B(n_319),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1037),
.Y(n_1096)
);

BUFx2_ASAP7_75t_SL g1097 ( 
.A(n_976),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_964),
.B(n_688),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_979),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_989),
.A2(n_986),
.B(n_1007),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1009),
.A2(n_200),
.B(n_316),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_977),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1033),
.A2(n_198),
.B(n_314),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1028),
.A2(n_197),
.B1(n_313),
.B2(n_310),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_1021),
.A2(n_1024),
.B(n_998),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1025),
.A2(n_1013),
.B(n_1011),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_972),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_992),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1078),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1089),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1039),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1038),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1091),
.B(n_995),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1077),
.A2(n_988),
.B1(n_985),
.B2(n_1019),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1049),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1089),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1084),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1085),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1058),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1057),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1087),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1040),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1070),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1107),
.A2(n_1032),
.B1(n_992),
.B2(n_1036),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1057),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1099),
.A2(n_992),
.B1(n_1002),
.B2(n_1029),
.Y(n_1126)
);

CKINVDCx11_ASAP7_75t_R g1127 ( 
.A(n_1050),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1040),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1044),
.A2(n_41),
.B(n_42),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1069),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1108),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1069),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1051),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1044),
.A2(n_318),
.B(n_69),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1043),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1059),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1102),
.A2(n_44),
.B1(n_70),
.B2(n_71),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1043),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_SL g1139 ( 
.A(n_1046),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1059),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1053),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1108),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1088),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1070),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1061),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1047),
.A2(n_97),
.B(n_99),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1079),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1067),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1104),
.A2(n_101),
.B1(n_106),
.B2(n_108),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_1067),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1079),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1079),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1046),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1064),
.A2(n_109),
.B(n_112),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1076),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1068),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1047),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1055),
.A2(n_113),
.B(n_115),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1076),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1102),
.A2(n_1066),
.B1(n_1097),
.B2(n_1105),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1066),
.A2(n_116),
.B1(n_118),
.B2(n_122),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1071),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1083),
.B(n_123),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1083),
.Y(n_1164)
);

CKINVDCx11_ASAP7_75t_R g1165 ( 
.A(n_1050),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1090),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1062),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_1066),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1096),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1041),
.B(n_1080),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1053),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1080),
.B(n_125),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1105),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1144),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_R g1175 ( 
.A(n_1115),
.B(n_1073),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1112),
.B(n_1082),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1113),
.B(n_1114),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1154),
.A2(n_1086),
.B1(n_1065),
.B2(n_1060),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1109),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1111),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1148),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1116),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1119),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1120),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1125),
.B(n_1167),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1117),
.Y(n_1186)
);

NAND2xp33_ASAP7_75t_R g1187 ( 
.A(n_1153),
.B(n_1073),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1121),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1114),
.B(n_1082),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1110),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1118),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1167),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1122),
.B(n_1098),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1127),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_R g1195 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1169),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1141),
.B(n_1054),
.Y(n_1197)
);

CKINVDCx11_ASAP7_75t_R g1198 ( 
.A(n_1127),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1162),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1148),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1128),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1162),
.Y(n_1202)
);

AO32x2_ASAP7_75t_L g1203 ( 
.A1(n_1143),
.A2(n_1131),
.A3(n_1129),
.B1(n_1160),
.B2(n_1124),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_R g1204 ( 
.A(n_1170),
.B(n_1093),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1119),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1171),
.B(n_1042),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1136),
.B(n_1063),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1136),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1137),
.B(n_1106),
.C(n_1072),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1146),
.A2(n_1094),
.B(n_1101),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1123),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1130),
.Y(n_1212)
);

NAND2x1_ASAP7_75t_L g1213 ( 
.A(n_1144),
.B(n_1056),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1139),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_R g1215 ( 
.A(n_1165),
.B(n_1042),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1123),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_R g1217 ( 
.A(n_1165),
.B(n_1042),
.Y(n_1217)
);

NAND3xp33_ASAP7_75t_L g1218 ( 
.A(n_1161),
.B(n_1092),
.C(n_1052),
.Y(n_1218)
);

NAND2xp33_ASAP7_75t_R g1219 ( 
.A(n_1159),
.B(n_1052),
.Y(n_1219)
);

AND2x2_ASAP7_75t_SL g1220 ( 
.A(n_1131),
.B(n_1081),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1145),
.B(n_1060),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1160),
.A2(n_1086),
.B1(n_1072),
.B2(n_1075),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1139),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1161),
.A2(n_1065),
.B1(n_1103),
.B2(n_1072),
.C1(n_1100),
.C2(n_1101),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1132),
.B(n_1075),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1149),
.A2(n_1100),
.B(n_1048),
.C(n_1103),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1168),
.B(n_1046),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1133),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1140),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1137),
.B(n_1052),
.C(n_1081),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1147),
.B(n_1074),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1151),
.B(n_1048),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1129),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1177),
.B(n_1152),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1198),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1233),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1212),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1221),
.B(n_1129),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1184),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1181),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1213),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1182),
.B(n_1126),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1208),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1192),
.B(n_1189),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1233),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1202),
.B(n_1166),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1180),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1186),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1201),
.B(n_1196),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1225),
.B(n_1126),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1191),
.B(n_1142),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1190),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1229),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1176),
.B(n_1163),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1205),
.B(n_1164),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1232),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1230),
.B(n_1173),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1179),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1188),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1231),
.B(n_1142),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1211),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1216),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1181),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1194),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1210),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1228),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1226),
.B(n_1135),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1207),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1199),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1220),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1183),
.B(n_1164),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1203),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1174),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1193),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1206),
.B(n_1164),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1219),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1222),
.B(n_1138),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1178),
.B(n_1157),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1209),
.B(n_1163),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1187),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1224),
.B(n_1156),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1174),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1200),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1200),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1185),
.B(n_1095),
.Y(n_1285)
);

INVx2_ASAP7_75t_R g1286 ( 
.A(n_1195),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1204),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1197),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1218),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1215),
.B(n_1095),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1247),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1236),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1236),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1245),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1287),
.B(n_1158),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1250),
.B(n_1134),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1288),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1286),
.B(n_1217),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1268),
.B(n_1227),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1245),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1238),
.B(n_1045),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1244),
.B(n_1214),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1248),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1237),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_1045),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1272),
.B(n_1164),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1253),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1257),
.B(n_1175),
.C(n_1155),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1243),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1276),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1274),
.B(n_1150),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1285),
.B(n_1223),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1280),
.A2(n_144),
.B1(n_146),
.B2(n_148),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1258),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1256),
.B(n_150),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1256),
.B(n_154),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1278),
.B(n_158),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1278),
.B(n_160),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1234),
.B(n_161),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1241),
.B(n_162),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_L g1321 ( 
.A(n_1266),
.B(n_166),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1269),
.B(n_167),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1242),
.B(n_169),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1286),
.B(n_178),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1277),
.B(n_180),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1277),
.B(n_1270),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1249),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1246),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1249),
.B(n_183),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1326),
.B(n_1285),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1326),
.B(n_1267),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1291),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1309),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1303),
.Y(n_1334)
);

AND2x2_ASAP7_75t_SL g1335 ( 
.A(n_1298),
.B(n_1279),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1328),
.B(n_1289),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1310),
.B(n_1270),
.Y(n_1337)
);

AND2x2_ASAP7_75t_SL g1338 ( 
.A(n_1295),
.B(n_1279),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1304),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1292),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1314),
.B(n_1260),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1307),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1312),
.B(n_1254),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1301),
.B(n_1305),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1327),
.B(n_1281),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1293),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1312),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1306),
.B(n_1265),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1306),
.B(n_1294),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1327),
.B(n_1249),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1300),
.B(n_1255),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1300),
.B(n_1290),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1336),
.B(n_1296),
.Y(n_1355)
);

AOI32xp33_ASAP7_75t_L g1356 ( 
.A1(n_1331),
.A2(n_1295),
.A3(n_1318),
.B1(n_1317),
.B2(n_1325),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1344),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1340),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1338),
.A2(n_1308),
.B(n_1257),
.C(n_1321),
.Y(n_1359)
);

NOR2x1_ASAP7_75t_R g1360 ( 
.A(n_1349),
.B(n_1264),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1343),
.B(n_1235),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1354),
.B(n_1331),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1349),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1330),
.B(n_1297),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1335),
.A2(n_1251),
.B1(n_1317),
.B2(n_1318),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1345),
.B(n_1297),
.Y(n_1366)
);

OA222x2_ASAP7_75t_L g1367 ( 
.A1(n_1337),
.A2(n_1341),
.B1(n_1347),
.B2(n_1324),
.C1(n_1353),
.C2(n_1339),
.Y(n_1367)
);

O2A1O1Ixp5_ASAP7_75t_R g1368 ( 
.A1(n_1352),
.A2(n_1299),
.B(n_1302),
.C(n_1311),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1340),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1332),
.Y(n_1370)
);

OAI211xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1334),
.A2(n_1322),
.B(n_1319),
.C(n_1271),
.Y(n_1371)
);

OAI211xp5_ASAP7_75t_L g1372 ( 
.A1(n_1368),
.A2(n_1359),
.B(n_1365),
.C(n_1356),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1370),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1358),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1369),
.Y(n_1375)
);

OAI31xp33_ASAP7_75t_L g1376 ( 
.A1(n_1361),
.A2(n_1320),
.A3(n_1313),
.B(n_1323),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1371),
.A2(n_1360),
.B(n_1355),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1366),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1355),
.B(n_1333),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1357),
.Y(n_1380)
);

AOI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1367),
.A2(n_1329),
.B(n_1323),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_SL g1382 ( 
.A(n_1372),
.B(n_1320),
.C(n_1342),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1373),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1380),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1378),
.B(n_1362),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1377),
.B(n_1239),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1381),
.A2(n_1363),
.B(n_1239),
.C(n_1346),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1374),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1375),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1376),
.B(n_1364),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1379),
.A2(n_1251),
.B(n_1315),
.Y(n_1391)
);

NOR3x1_ASAP7_75t_L g1392 ( 
.A(n_1382),
.B(n_1275),
.C(n_1284),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1383),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1388),
.B(n_1351),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1387),
.B(n_1391),
.Y(n_1396)
);

OA22x2_ASAP7_75t_L g1397 ( 
.A1(n_1390),
.A2(n_1351),
.B1(n_1348),
.B2(n_1350),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1396),
.A2(n_1389),
.B(n_1384),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1393),
.B(n_1316),
.C(n_1259),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1394),
.B(n_1397),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1395),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1401),
.Y(n_1402)
);

OAI222xp33_ASAP7_75t_L g1403 ( 
.A1(n_1400),
.A2(n_1392),
.B1(n_1316),
.B2(n_1283),
.C1(n_1241),
.C2(n_1282),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1398),
.A2(n_1262),
.B(n_1261),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1399),
.A2(n_1252),
.B1(n_1263),
.B2(n_1240),
.C(n_1273),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1402),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1404),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_L g1408 ( 
.A(n_1403),
.B(n_1263),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1405),
.Y(n_1409)
);

AND3x2_ASAP7_75t_L g1410 ( 
.A(n_1406),
.B(n_184),
.C(n_193),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1409),
.A2(n_1240),
.B1(n_201),
.B2(n_207),
.C(n_208),
.Y(n_1411)
);

NAND2x1_ASAP7_75t_SL g1412 ( 
.A(n_1408),
.B(n_196),
.Y(n_1412)
);

OR3x2_ASAP7_75t_L g1413 ( 
.A(n_1407),
.B(n_211),
.C(n_214),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1412),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1413),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1410),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1411),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1416),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1414),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1415),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1420),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1418),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1419),
.A2(n_1417),
.B1(n_223),
.B2(n_228),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1422),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1421),
.B(n_218),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1423),
.A2(n_236),
.B(n_242),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1424),
.A2(n_250),
.B1(n_253),
.B2(n_255),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1426),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1425),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1428),
.A2(n_1427),
.B1(n_263),
.B2(n_268),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1429),
.A2(n_262),
.B(n_269),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1430),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1431),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1432),
.A2(n_295),
.B1(n_296),
.B2(n_300),
.C(n_301),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1434),
.A2(n_1433),
.B1(n_304),
.B2(n_307),
.Y(n_1435)
);


endmodule