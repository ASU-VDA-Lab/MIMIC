module fake_ariane_1281_n_1708 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1708);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1708;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_36),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_18),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_59),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_27),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_20),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_20),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_58),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_21),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_22),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_100),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_66),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_56),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_24),
.Y(n_191)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_121),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_25),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_79),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_67),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_94),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_19),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_143),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_49),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_84),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_107),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_60),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_72),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_69),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_44),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_31),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_28),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_77),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_139),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_105),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_65),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_54),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_4),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_64),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_15),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_151),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_21),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_110),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_52),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_70),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_97),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_9),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_119),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_31),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_148),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_124),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_43),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_53),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_127),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_39),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_108),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_38),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_113),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_99),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_114),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_131),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_96),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_12),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_106),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_109),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_86),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_17),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_43),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_51),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_154),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_152),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_153),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_30),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_11),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_41),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_10),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_145),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_118),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_78),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_28),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_176),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_176),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_193),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_164),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_239),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_164),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_176),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_176),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_265),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_205),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_211),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_275),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_234),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_158),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_183),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_236),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_163),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_205),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_170),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_276),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_189),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_237),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_218),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_250),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_222),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_223),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_224),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_158),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_241),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_242),
.Y(n_367)
);

INVx4_ASAP7_75t_SL g368 ( 
.A(n_294),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_159),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_225),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_227),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_159),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_165),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_245),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_243),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_256),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_262),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_248),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_293),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_304),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_249),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_314),
.A2(n_291),
.B1(n_292),
.B2(n_284),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_316),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_247),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_371),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_342),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_R g403 ( 
.A(n_365),
.B(n_165),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_315),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_317),
.B(n_251),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_339),
.B(n_208),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_327),
.B(n_300),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_340),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_343),
.B(n_266),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_344),
.B(n_346),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_280),
.B1(n_191),
.B2(n_308),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_341),
.B(n_306),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_326),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_331),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_359),
.B(n_163),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_330),
.A2(n_179),
.B1(n_166),
.B2(n_308),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_352),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_355),
.B(n_157),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_366),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_383),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_389),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_367),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

AND3x2_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_369),
.C(n_336),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_359),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_375),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_378),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_373),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_423),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_167),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

AND3x2_ASAP7_75t_L g480 ( 
.A(n_391),
.B(n_345),
.C(n_221),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_401),
.B(n_361),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_361),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_392),
.B(n_171),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_368),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_405),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_368),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_401),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_424),
.B(n_156),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_362),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_410),
.Y(n_506)
);

INVx8_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_388),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_405),
.A2(n_310),
.B1(n_186),
.B2(n_172),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_368),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_400),
.B(n_156),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_415),
.B(n_362),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_402),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_422),
.B(n_363),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_409),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_415),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_400),
.B(n_161),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_405),
.A2(n_197),
.B1(n_186),
.B2(n_172),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_380),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_413),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_387),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_417),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_404),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_395),
.B(n_380),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_387),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_432),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_387),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_422),
.B(n_363),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_382),
.B(n_368),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_400),
.B(n_161),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_382),
.B(n_370),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_382),
.B(n_370),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_386),
.B(n_171),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_162),
.Y(n_558)
);

BUFx6f_ASAP7_75t_SL g559 ( 
.A(n_420),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_404),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_404),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_395),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_419),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_404),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_408),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_408),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_408),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_418),
.B(n_162),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_402),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_408),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_408),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_419),
.Y(n_577)
);

CKINVDCx6p67_ASAP7_75t_R g578 ( 
.A(n_393),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_420),
.B(n_374),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_406),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_419),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_433),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_420),
.B(n_374),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_418),
.B(n_168),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_420),
.B(n_376),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_433),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

AO21x2_ASAP7_75t_L g589 ( 
.A1(n_416),
.A2(n_178),
.B(n_169),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_436),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_436),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_447),
.B(n_444),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_411),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_484),
.B(n_444),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_475),
.B(n_411),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_527),
.B(n_471),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_527),
.B(n_393),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_477),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_494),
.B(n_430),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_494),
.B(n_425),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_478),
.B(n_411),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_478),
.B(n_416),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_536),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_565),
.A2(n_437),
.B(n_428),
.C(n_429),
.Y(n_607)
);

AND2x2_ASAP7_75t_SL g608 ( 
.A(n_558),
.B(n_181),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_478),
.B(n_427),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_477),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_499),
.B(n_427),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_478),
.A2(n_403),
.B1(n_421),
.B2(n_438),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_586),
.A2(n_438),
.B(n_437),
.C(n_429),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_494),
.B(n_439),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_592),
.B(n_428),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_478),
.B(n_445),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_478),
.B(n_446),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_531),
.B(n_168),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_531),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_478),
.B(n_446),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_531),
.B(n_173),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_544),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_531),
.B(n_173),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_472),
.B(n_528),
.C(n_520),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_499),
.B(n_439),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_477),
.A2(n_446),
.B1(n_386),
.B2(n_197),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_449),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_521),
.B(n_174),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_523),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_521),
.B(n_160),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_524),
.B(n_174),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_450),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_549),
.B(n_253),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_403),
.C(n_231),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_507),
.B(n_254),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_507),
.A2(n_559),
.B1(n_547),
.B2(n_504),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_532),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_507),
.B(n_175),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_507),
.B(n_175),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_546),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_450),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_451),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_451),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_589),
.A2(n_186),
.B1(n_235),
.B2(n_197),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_509),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_559),
.B(n_259),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_573),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_509),
.B(n_376),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_579),
.B(n_177),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_584),
.B(n_177),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_541),
.B(n_180),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_559),
.B(n_191),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_542),
.B(n_182),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_592),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_589),
.B(n_481),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_465),
.B(n_187),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_452),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_187),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_452),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_470),
.B(n_188),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_580),
.B(n_231),
.C(n_298),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_532),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_454),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_458),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_581),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_545),
.B(n_553),
.Y(n_670)
);

OAI221xp5_ASAP7_75t_L g671 ( 
.A1(n_517),
.A2(n_270),
.B1(n_301),
.B2(n_288),
.C(n_303),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_532),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_481),
.B(n_188),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_454),
.A2(n_377),
.B(n_379),
.C(n_329),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_532),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_572),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_585),
.B(n_270),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_460),
.A2(n_379),
.B(n_329),
.C(n_338),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_545),
.A2(n_233),
.B(n_228),
.C(n_216),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_553),
.B(n_273),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_467),
.B(n_431),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_467),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_555),
.B(n_273),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_581),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_581),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_550),
.B(n_551),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_460),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_543),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_594),
.B(n_184),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_467),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_555),
.B(n_271),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_467),
.B(n_431),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_564),
.B(n_426),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_SL g694 ( 
.A(n_543),
.B(n_285),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_529),
.B(n_285),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_487),
.B(n_298),
.C(n_288),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_594),
.B(n_566),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_594),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_505),
.A2(n_274),
.B1(n_277),
.B2(n_278),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

AOI221xp5_ASAP7_75t_L g701 ( 
.A1(n_557),
.A2(n_301),
.B1(n_303),
.B2(n_305),
.C(n_337),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_448),
.B(n_305),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_566),
.B(n_271),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_491),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_468),
.B(n_469),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_491),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_577),
.B(n_274),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_448),
.B(n_277),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_493),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_577),
.B(n_279),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_458),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_505),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_493),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_582),
.B(n_281),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_468),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_469),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_483),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_582),
.B(n_290),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_583),
.B(n_290),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_295),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_458),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_483),
.A2(n_525),
.B(n_533),
.C(n_501),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_465),
.B(n_295),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_578),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_578),
.B(n_426),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_498),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_490),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_590),
.B(n_453),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_465),
.B(n_309),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_505),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_590),
.B(n_309),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_490),
.Y(n_732)
);

INVx8_ASAP7_75t_L g733 ( 
.A(n_465),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_448),
.B(n_185),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_465),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_476),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_476),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_453),
.B(n_199),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_476),
.B(n_190),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_557),
.B(n_464),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_496),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_496),
.A2(n_235),
.B1(n_163),
.B2(n_172),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_457),
.B(n_201),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_455),
.B(n_194),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_457),
.B(n_202),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_476),
.B(n_196),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_455),
.B(n_215),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_459),
.B(n_203),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_502),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_459),
.B(n_204),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_500),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_461),
.B(n_206),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_455),
.B(n_252),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_587),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_476),
.B(n_255),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_479),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_502),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_479),
.B(n_263),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_500),
.A2(n_235),
.B1(n_332),
.B2(n_338),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_501),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_606),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_630),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_647),
.B(n_480),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_611),
.B(n_587),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_608),
.A2(n_593),
.B1(n_591),
.B2(n_588),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_628),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_461),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_611),
.B(n_588),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_724),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_667),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_633),
.B(n_591),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_643),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_639),
.B(n_463),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_608),
.B(n_479),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_644),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_619),
.B(n_479),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_660),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_619),
.B(n_479),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_682),
.B(n_511),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_662),
.B(n_666),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_687),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_SL g784 ( 
.A1(n_627),
.A2(n_695),
.B1(n_692),
.B2(n_681),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_693),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_672),
.B(n_650),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_SL g787 ( 
.A(n_711),
.B(n_511),
.C(n_539),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_715),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_682),
.B(n_512),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_725),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_690),
.B(n_512),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_627),
.A2(n_593),
.B1(n_503),
.B2(n_506),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_636),
.B(n_514),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_690),
.B(n_514),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_717),
.B(n_522),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_623),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_SL g800 ( 
.A1(n_695),
.A2(n_335),
.B1(n_334),
.B2(n_332),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_603),
.A2(n_675),
.B1(n_665),
.B2(n_632),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_598),
.B(n_488),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_727),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_732),
.B(n_522),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_735),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_665),
.B(n_488),
.Y(n_807)
);

BUFx8_ASAP7_75t_L g808 ( 
.A(n_681),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_741),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_638),
.B(n_489),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_692),
.Y(n_811)
);

AO22x1_ASAP7_75t_L g812 ( 
.A1(n_730),
.A2(n_518),
.B1(n_497),
.B2(n_335),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_735),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_688),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_712),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_751),
.B(n_525),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_740),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_675),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_737),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_760),
.B(n_658),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_686),
.B(n_533),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_634),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_596),
.B(n_535),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_700),
.B(n_535),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_637),
.A2(n_609),
.B1(n_605),
.B2(n_596),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_700),
.B(n_538),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_722),
.B(n_705),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_642),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_614),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_601),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_712),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_595),
.B(n_538),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_637),
.B(n_488),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_599),
.B(n_463),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_610),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_620),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_699),
.B(n_640),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_684),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_625),
.B(n_539),
.Y(n_839)
);

BUFx4f_ASAP7_75t_L g840 ( 
.A(n_689),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_597),
.B(n_607),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_652),
.B(n_466),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_646),
.A2(n_506),
.B1(n_513),
.B2(n_508),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_646),
.A2(n_503),
.B1(n_513),
.B2(n_508),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_694),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_685),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_641),
.B(n_655),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_SL g848 ( 
.A(n_677),
.B(n_296),
.C(n_272),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_602),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_631),
.B(n_334),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_600),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_615),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_728),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_663),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_604),
.B(n_466),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_668),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_704),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_655),
.Y(n_859)
);

NOR2x2_ASAP7_75t_L g860 ( 
.A(n_701),
.B(n_473),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_626),
.B(n_473),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_664),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_735),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_625),
.B(n_482),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_673),
.B(n_337),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_612),
.B(n_488),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_652),
.B(n_482),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_677),
.B(n_485),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_629),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_709),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_726),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_657),
.B(n_492),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_657),
.B(n_648),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_648),
.B(n_492),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_652),
.B(n_485),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_735),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_749),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_757),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_635),
.A2(n_486),
.B1(n_510),
.B2(n_516),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_689),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_669),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_669),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_754),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_697),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_SL g887 ( 
.A(n_696),
.B(n_229),
.C(n_207),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_618),
.B(n_492),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_618),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_622),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_622),
.B(n_492),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_742),
.B(n_515),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_624),
.B(n_492),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_624),
.B(n_486),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_652),
.B(n_526),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_652),
.B(n_526),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_635),
.B(n_456),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_742),
.A2(n_510),
.B1(n_516),
.B2(n_474),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_736),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_652),
.B(n_495),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_613),
.B(n_456),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_736),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_736),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_702),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_661),
.A2(n_671),
.B1(n_759),
.B2(n_616),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_737),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_756),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_678),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_756),
.B(n_456),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_680),
.B(n_474),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_676),
.B(n_474),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_670),
.A2(n_515),
.B(n_516),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_617),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_654),
.B(n_519),
.C(n_495),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_621),
.B(n_510),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_680),
.B(n_571),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_651),
.B(n_653),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_683),
.B(n_571),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_702),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_683),
.B(n_571),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_674),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_708),
.A2(n_519),
.B1(n_495),
.B2(n_515),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_759),
.B(n_560),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_656),
.B(n_495),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_739),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_708),
.A2(n_519),
.B1(n_495),
.B2(n_574),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_703),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_691),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_707),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_734),
.B(n_560),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_734),
.B(n_519),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_710),
.B(n_519),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_714),
.B(n_552),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_718),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_744),
.B(n_561),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_719),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_561),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_739),
.B(n_562),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_720),
.B(n_552),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_731),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_747),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_766),
.Y(n_942)
);

NAND2x2_ASAP7_75t_L g943 ( 
.A(n_763),
.B(n_738),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_821),
.B(n_747),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_814),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_770),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_825),
.A2(n_753),
.B(n_679),
.C(n_748),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_761),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_821),
.A2(n_753),
.B1(n_659),
.B2(n_750),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_772),
.Y(n_950)
);

AO221x1_ASAP7_75t_L g951 ( 
.A1(n_784),
.A2(n_307),
.B1(n_282),
.B2(n_287),
.C(n_297),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_823),
.A2(n_659),
.B(n_723),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_R g953 ( 
.A(n_792),
.B(n_743),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_904),
.A2(n_745),
.B(n_752),
.C(n_575),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_808),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_859),
.B(n_729),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_769),
.Y(n_957)
);

OAI22x1_ASAP7_75t_L g958 ( 
.A1(n_811),
.A2(n_758),
.B1(n_755),
.B2(n_746),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_776),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_823),
.A2(n_576),
.B(n_540),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_848),
.A2(n_758),
.B(n_755),
.C(n_746),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_802),
.A2(n_563),
.B(n_575),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_798),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_832),
.A2(n_576),
.B(n_540),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_762),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_774),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_840),
.B(n_919),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_762),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_820),
.B(n_562),
.Y(n_969)
);

OAI22x1_ASAP7_75t_L g970 ( 
.A1(n_889),
.A2(n_299),
.B1(n_302),
.B2(n_569),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_789),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_789),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_799),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_822),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_824),
.B(n_563),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_824),
.B(n_568),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_828),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_857),
.Y(n_978)
);

BUFx12f_ASAP7_75t_L g979 ( 
.A(n_808),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_826),
.B(n_568),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_895),
.A2(n_574),
.B(n_570),
.Y(n_981)
);

AOI221xp5_ASAP7_75t_L g982 ( 
.A1(n_848),
.A2(n_192),
.B1(n_569),
.B2(n_570),
.C(n_238),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_895),
.A2(n_896),
.B(n_841),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_785),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_896),
.A2(n_530),
.B(n_556),
.Y(n_985)
);

CKINVDCx10_ASAP7_75t_R g986 ( 
.A(n_845),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_778),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_861),
.A2(n_567),
.B(n_552),
.C(n_548),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_799),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_841),
.A2(n_556),
.B(n_554),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_567),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_837),
.A2(n_567),
.B(n_552),
.C(n_554),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_904),
.A2(n_0),
.B(n_2),
.C(n_5),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_SL g994 ( 
.A1(n_928),
.A2(n_567),
.B(n_552),
.C(n_7),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_764),
.A2(n_556),
.B(n_554),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_818),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_779),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_847),
.B(n_209),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_927),
.B(n_212),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_797),
.A2(n_213),
.B1(n_214),
.B2(n_217),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_854),
.B(n_537),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_764),
.A2(n_537),
.B(n_534),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_840),
.B(n_246),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_768),
.A2(n_827),
.B(n_842),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_SL g1005 ( 
.A1(n_800),
.A2(n_219),
.B1(n_220),
.B2(n_226),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_882),
.B(n_537),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_781),
.B(n_257),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_768),
.A2(n_534),
.B(n_530),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_781),
.B(n_264),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_783),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_801),
.A2(n_230),
.B1(n_232),
.B2(n_240),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_917),
.A2(n_0),
.B(n_6),
.C(n_8),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_787),
.B(n_244),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_790),
.B(n_268),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_851),
.B(n_6),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_817),
.B(n_8),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_871),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_788),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_790),
.B(n_385),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_787),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_793),
.B(n_534),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_791),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_827),
.A2(n_530),
.B(n_385),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_793),
.B(n_385),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_929),
.A2(n_385),
.B(n_14),
.C(n_15),
.Y(n_1025)
);

AOI33xp33_ASAP7_75t_L g1026 ( 
.A1(n_936),
.A2(n_13),
.A3(n_16),
.B1(n_22),
.B2(n_23),
.B3(n_24),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_842),
.A2(n_385),
.B(n_442),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_797),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_803),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_829),
.B(n_29),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_805),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_852),
.A2(n_385),
.B1(n_42),
.B2(n_45),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_941),
.B(n_37),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_853),
.B(n_385),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_796),
.B(n_385),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_940),
.A2(n_42),
.B(n_45),
.C(n_48),
.Y(n_1036)
);

NAND3x1_ASAP7_75t_L g1037 ( 
.A(n_767),
.B(n_73),
.C(n_76),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_941),
.A2(n_80),
.B(n_82),
.C(n_88),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_886),
.B(n_95),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_805),
.A2(n_101),
.B1(n_117),
.B2(n_120),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_SL g1041 ( 
.A1(n_892),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_1041)
);

CKINVDCx6p67_ASAP7_75t_R g1042 ( 
.A(n_862),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_879),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_809),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_858),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_816),
.A2(n_138),
.B1(n_141),
.B2(n_147),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_855),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_816),
.A2(n_782),
.B1(n_839),
.B2(n_921),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_863),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_866),
.B(n_885),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_868),
.A2(n_877),
.B(n_937),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_860),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_872),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_799),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_782),
.B(n_839),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_804),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_928),
.A2(n_911),
.B(n_918),
.C(n_910),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_934),
.B(n_869),
.Y(n_1059)
);

CKINVDCx6p67_ASAP7_75t_R g1060 ( 
.A(n_864),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_901),
.A2(n_930),
.B(n_935),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_R g1062 ( 
.A(n_804),
.B(n_899),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_795),
.A2(n_890),
.B(n_834),
.C(n_865),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_870),
.A2(n_880),
.B1(n_850),
.B2(n_905),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_838),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_875),
.B(n_796),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_804),
.B(n_899),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_902),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_864),
.B(n_878),
.Y(n_1069)
);

OAI321xp33_ASAP7_75t_L g1070 ( 
.A1(n_908),
.A2(n_775),
.A3(n_910),
.B1(n_916),
.B2(n_918),
.C(n_920),
.Y(n_1070)
);

CKINVDCx11_ASAP7_75t_R g1071 ( 
.A(n_806),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_846),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_849),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_815),
.B(n_831),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_771),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_830),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_868),
.A2(n_877),
.B(n_937),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_865),
.A2(n_897),
.B(n_773),
.C(n_916),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_930),
.A2(n_935),
.B(n_912),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_771),
.B(n_913),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1071),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_944),
.A2(n_983),
.B(n_1051),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1079),
.A2(n_912),
.B(n_901),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1048),
.A2(n_920),
.B1(n_887),
.B2(n_881),
.Y(n_1084)
);

CKINVDCx8_ASAP7_75t_R g1085 ( 
.A(n_986),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_900),
.B(n_924),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1048),
.A2(n_867),
.B(n_922),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1004),
.A2(n_939),
.B(n_932),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1056),
.B(n_835),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_1028),
.A2(n_925),
.A3(n_907),
.B1(n_887),
.B2(n_812),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1060),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_1033),
.A2(n_894),
.B(n_909),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_988),
.A2(n_923),
.A3(n_925),
.B(n_836),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1052),
.B(n_786),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1061),
.A2(n_914),
.B(n_833),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_942),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_945),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_962),
.A2(n_981),
.B(n_992),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_SL g1099 ( 
.A(n_1041),
.B(n_931),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1056),
.B(n_883),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_965),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_955),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_996),
.B(n_884),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_984),
.B(n_898),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1061),
.A2(n_1023),
.B(n_990),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_947),
.A2(n_926),
.B(n_931),
.Y(n_1106)
);

OAI22x1_ASAP7_75t_L g1107 ( 
.A1(n_1032),
.A2(n_876),
.B1(n_893),
.B2(n_891),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_952),
.A2(n_888),
.B(n_874),
.Y(n_1108)
);

NOR4xp25_ASAP7_75t_L g1109 ( 
.A(n_1028),
.B(n_807),
.C(n_923),
.D(n_844),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_946),
.B(n_903),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_971),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1070),
.A2(n_931),
.B(n_915),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1047),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_998),
.A2(n_915),
.B(n_906),
.C(n_938),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1016),
.B(n_938),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_1058),
.A2(n_777),
.B(n_780),
.C(n_819),
.Y(n_1116)
);

NAND3x1_ASAP7_75t_L g1117 ( 
.A(n_1026),
.B(n_819),
.C(n_933),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_964),
.A2(n_843),
.B(n_765),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_960),
.A2(n_864),
.B(n_878),
.Y(n_1119)
);

AO32x2_ASAP7_75t_L g1120 ( 
.A1(n_1031),
.A2(n_810),
.A3(n_931),
.B1(n_794),
.B2(n_856),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_949),
.A2(n_878),
.B(n_813),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1078),
.A2(n_810),
.A3(n_856),
.B(n_913),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1021),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_949),
.A2(n_806),
.B(n_813),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1006),
.B(n_909),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1070),
.A2(n_806),
.B(n_913),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_985),
.A2(n_969),
.B(n_1027),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_969),
.A2(n_810),
.B(n_856),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1021),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_958),
.A2(n_856),
.A3(n_1039),
.B(n_1075),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1039),
.A2(n_1080),
.B(n_1008),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1015),
.A2(n_1031),
.B1(n_1030),
.B2(n_1044),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_979),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_966),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_951),
.A2(n_1005),
.B1(n_1011),
.B2(n_1066),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_995),
.A2(n_1002),
.B(n_1038),
.Y(n_1136)
);

BUFx8_ASAP7_75t_L g1137 ( 
.A(n_971),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1063),
.A2(n_1001),
.B(n_961),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_SL g1139 ( 
.A(n_971),
.B(n_1055),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_SL g1140 ( 
.A1(n_1020),
.A2(n_993),
.B(n_991),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_SL g1141 ( 
.A1(n_1040),
.A2(n_1046),
.B(n_1073),
.C(n_1072),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_968),
.Y(n_1142)
);

OA21x2_ASAP7_75t_L g1143 ( 
.A1(n_1001),
.A2(n_982),
.B(n_1036),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1037),
.A2(n_1040),
.B(n_1046),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1059),
.B(n_1050),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_1049),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_970),
.A2(n_1053),
.A3(n_948),
.B(n_1017),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1076),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_999),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_954),
.A2(n_994),
.B(n_1069),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1012),
.A2(n_1064),
.B(n_1059),
.C(n_1010),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_963),
.A2(n_977),
.A3(n_974),
.B(n_978),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1000),
.A2(n_1042),
.B1(n_967),
.B2(n_1009),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1000),
.A2(n_980),
.B1(n_976),
.B2(n_975),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_953),
.Y(n_1155)
);

AOI211x1_ASAP7_75t_L g1156 ( 
.A1(n_950),
.A2(n_1022),
.B(n_959),
.C(n_1018),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1034),
.A2(n_1065),
.B(n_1029),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_987),
.A2(n_997),
.B(n_1019),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1068),
.B(n_1043),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1055),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1007),
.B(n_1014),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1024),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1062),
.Y(n_1163)
);

AOI221x1_ASAP7_75t_L g1164 ( 
.A1(n_972),
.A2(n_973),
.B1(n_989),
.B2(n_1024),
.C(n_1035),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_1035),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_943),
.A2(n_1003),
.B1(n_1006),
.B2(n_1067),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_973),
.B(n_989),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1074),
.Y(n_1168)
);

AO32x2_ASAP7_75t_L g1169 ( 
.A1(n_1057),
.A2(n_1048),
.A3(n_1031),
.B1(n_1028),
.B2(n_784),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1013),
.A2(n_944),
.B(n_904),
.C(n_1058),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1006),
.B(n_688),
.Y(n_1171)
);

AND2x6_ASAP7_75t_SL g1172 ( 
.A(n_956),
.B(n_467),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1054),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_944),
.A2(n_983),
.B(n_823),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1052),
.B(n_565),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1056),
.B(n_688),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1056),
.B(n_688),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1071),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_946),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1048),
.A2(n_848),
.B1(n_608),
.B2(n_565),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1056),
.B(n_688),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1079),
.A2(n_962),
.B(n_983),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1052),
.B(n_647),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_944),
.A2(n_983),
.B(n_823),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1048),
.A2(n_447),
.B(n_608),
.C(n_475),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1079),
.A2(n_1051),
.A3(n_1077),
.B(n_1048),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_688),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1048),
.A2(n_1078),
.B(n_944),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_955),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1056),
.B(n_688),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1079),
.A2(n_962),
.B(n_983),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1079),
.A2(n_962),
.B(n_983),
.Y(n_1192)
);

NAND2x1_ASAP7_75t_L g1193 ( 
.A(n_1075),
.B(n_819),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_996),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_962),
.B(n_983),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_951),
.A2(n_565),
.B1(n_784),
.B2(n_608),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1056),
.B(n_688),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1048),
.A2(n_447),
.B(n_608),
.C(n_475),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_996),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1048),
.A2(n_447),
.B(n_608),
.C(n_475),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1048),
.A2(n_944),
.B1(n_608),
.B2(n_1056),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1048),
.A2(n_447),
.B(n_608),
.C(n_475),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_957),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_944),
.A2(n_983),
.B(n_823),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1054),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_942),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1048),
.B(n_840),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1048),
.A2(n_848),
.B1(n_608),
.B2(n_565),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1052),
.B(n_647),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1079),
.A2(n_1051),
.A3(n_1077),
.B(n_1048),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1180),
.A2(n_1208),
.B1(n_1196),
.B2(n_1201),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1203),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1201),
.A2(n_1082),
.A3(n_1084),
.B(n_1174),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1198),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1202),
.A2(n_1180),
.B1(n_1208),
.B2(n_1135),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1132),
.A2(n_1188),
.B1(n_1109),
.B2(n_1149),
.C(n_1084),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1182),
.A2(n_1192),
.B(n_1191),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1144),
.A2(n_1099),
.B(n_1106),
.C(n_1132),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1195),
.A2(n_1105),
.B(n_1098),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1135),
.A2(n_1153),
.B1(n_1101),
.B2(n_1117),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1085),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1170),
.A2(n_1151),
.B(n_1207),
.C(n_1106),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1127),
.A2(n_1083),
.B(n_1136),
.Y(n_1224)
);

OAI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1153),
.A2(n_1099),
.B1(n_1109),
.B2(n_1087),
.C(n_1161),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1133),
.B(n_1189),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1125),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1088),
.A2(n_1086),
.B(n_1131),
.Y(n_1228)
);

BUFx4_ASAP7_75t_R g1229 ( 
.A(n_1134),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_1204),
.B(n_1184),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1141),
.A2(n_1126),
.B(n_1095),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1175),
.A2(n_1104),
.B1(n_1115),
.B2(n_1145),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1124),
.A2(n_1121),
.B(n_1138),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1112),
.A2(n_1169),
.B(n_1158),
.C(n_1114),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1173),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1179),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1112),
.A2(n_1150),
.B(n_1128),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1123),
.B(n_1129),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1093),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1118),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1143),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_1157),
.B(n_1100),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1089),
.A2(n_1206),
.B(n_1154),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1107),
.A2(n_1146),
.B(n_1143),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1102),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1103),
.B(n_1168),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1102),
.B(n_1183),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1093),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1123),
.B(n_1129),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1177),
.A2(n_1190),
.B(n_1181),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1093),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1187),
.B(n_1197),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1092),
.A2(n_1193),
.B(n_1146),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1186),
.A2(n_1210),
.B(n_1164),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1166),
.A2(n_1199),
.B1(n_1194),
.B2(n_1097),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1139),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_SL g1258 ( 
.A1(n_1171),
.A2(n_1167),
.B(n_1166),
.C(n_1110),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1156),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1162),
.B(n_1091),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1159),
.B(n_1205),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1137),
.Y(n_1262)
);

BUFx8_ASAP7_75t_L g1263 ( 
.A(n_1081),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1186),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1091),
.B(n_1160),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1137),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1091),
.B(n_1111),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1081),
.B(n_1178),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1186),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1081),
.B(n_1178),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1209),
.A2(n_1155),
.B(n_1094),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1120),
.A2(n_1210),
.B(n_1130),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1169),
.A2(n_1120),
.B(n_1090),
.C(n_1163),
.Y(n_1273)
);

BUFx4f_ASAP7_75t_L g1274 ( 
.A(n_1178),
.Y(n_1274)
);

AND2x6_ASAP7_75t_SL g1275 ( 
.A(n_1102),
.B(n_1113),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1210),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1152),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1147),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1120),
.A2(n_1130),
.B(n_1169),
.Y(n_1279)
);

BUFx2_ASAP7_75t_SL g1280 ( 
.A(n_1111),
.Y(n_1280)
);

INVx4_ASAP7_75t_SL g1281 ( 
.A(n_1122),
.Y(n_1281)
);

AOI222xp33_ASAP7_75t_L g1282 ( 
.A1(n_1172),
.A2(n_784),
.B1(n_565),
.B2(n_627),
.C1(n_557),
.C2(n_701),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1130),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1122),
.A2(n_1090),
.B(n_1172),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1090),
.B(n_1147),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1198),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1145),
.B(n_1194),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1137),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1145),
.B(n_1176),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1111),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_1133),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1145),
.B(n_1194),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1185),
.B(n_1198),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1180),
.A2(n_784),
.B1(n_951),
.B2(n_1208),
.Y(n_1296)
);

NOR2x1_ASAP7_75t_SL g1297 ( 
.A(n_1207),
.B(n_1048),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1185),
.A2(n_1198),
.B(n_1202),
.C(n_1200),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1148),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_784),
.B1(n_951),
.B2(n_1208),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1096),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1145),
.B(n_1176),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1198),
.Y(n_1304)
);

INVx8_ASAP7_75t_L g1305 ( 
.A(n_1133),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1185),
.A2(n_1200),
.B1(n_1202),
.B2(n_1198),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1185),
.A2(n_1198),
.B(n_1202),
.C(n_1200),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1145),
.B(n_1176),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1311)
);

INVx3_ASAP7_75t_SL g1312 ( 
.A(n_1179),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1185),
.B(n_1200),
.C(n_1198),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1098),
.A2(n_1191),
.B(n_1182),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1145),
.B(n_1194),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1096),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1085),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1198),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1096),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1202),
.C(n_1198),
.Y(n_1321)
);

NAND2x1_ASAP7_75t_L g1322 ( 
.A(n_1188),
.B(n_1138),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1182),
.A2(n_1192),
.B(n_1191),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1149),
.B(n_565),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1264),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1211),
.B(n_1237),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1231),
.A2(n_1286),
.B(n_1319),
.C(n_1215),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_L g1329 ( 
.A1(n_1294),
.A2(n_1306),
.B(n_1304),
.C(n_1321),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1264),
.A2(n_1276),
.B(n_1269),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1211),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1316),
.B(n_1247),
.Y(n_1332)
);

O2A1O1Ixp5_ASAP7_75t_L g1333 ( 
.A1(n_1294),
.A2(n_1304),
.B(n_1321),
.C(n_1322),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1267),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1253),
.B(n_1289),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1232),
.B(n_1237),
.Y(n_1336)
);

AOI31xp33_ASAP7_75t_L g1337 ( 
.A1(n_1217),
.A2(n_1296),
.A3(n_1301),
.B(n_1216),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1242),
.A2(n_1224),
.B(n_1255),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1217),
.A2(n_1223),
.B(n_1225),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1232),
.B(n_1300),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1303),
.B(n_1310),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1262),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1314),
.A2(n_1219),
.B(n_1233),
.C(n_1255),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_L g1344 ( 
.A(n_1246),
.B(n_1288),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1227),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1262),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1240),
.A2(n_1249),
.B(n_1252),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1296),
.A2(n_1301),
.B1(n_1212),
.B2(n_1225),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1308),
.A2(n_1221),
.B(n_1219),
.C(n_1298),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1242),
.A2(n_1245),
.B(n_1228),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1222),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1308),
.A2(n_1298),
.B(n_1230),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1251),
.B(n_1302),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1300),
.B(n_1309),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1317),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1240),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1223),
.A2(n_1282),
.B(n_1324),
.C(n_1256),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1320),
.B(n_1261),
.Y(n_1358)
);

AND2x2_ASAP7_75t_SL g1359 ( 
.A(n_1279),
.B(n_1212),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1234),
.A2(n_1324),
.B1(n_1273),
.B2(n_1262),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1227),
.B(n_1213),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1244),
.B(n_1239),
.Y(n_1362)
);

O2A1O1Ixp5_ASAP7_75t_L g1363 ( 
.A1(n_1273),
.A2(n_1234),
.B(n_1257),
.C(n_1284),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1318),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1259),
.B(n_1285),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1250),
.B(n_1265),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1244),
.B(n_1250),
.Y(n_1367)
);

BUFx8_ASAP7_75t_SL g1368 ( 
.A(n_1274),
.Y(n_1368)
);

BUFx2_ASAP7_75t_SL g1369 ( 
.A(n_1236),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1268),
.B(n_1270),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_SL g1371 ( 
.A(n_1263),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1257),
.A2(n_1274),
.B1(n_1271),
.B2(n_1266),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1268),
.B(n_1270),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1297),
.A2(n_1230),
.B(n_1260),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1284),
.A2(n_1312),
.B1(n_1292),
.B2(n_1229),
.Y(n_1375)
);

O2A1O1Ixp5_ASAP7_75t_L g1376 ( 
.A1(n_1291),
.A2(n_1278),
.B(n_1283),
.C(n_1260),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1243),
.A2(n_1241),
.B(n_1238),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1291),
.B(n_1280),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1218),
.A2(n_1323),
.B(n_1258),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1312),
.A2(n_1305),
.B1(n_1272),
.B2(n_1248),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1258),
.A2(n_1226),
.B(n_1272),
.C(n_1220),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1290),
.A2(n_1315),
.B(n_1313),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1220),
.A2(n_1235),
.B(n_1299),
.C(n_1214),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1214),
.A2(n_1275),
.B(n_1277),
.C(n_1305),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1305),
.A2(n_1214),
.B1(n_1263),
.B2(n_1254),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1295),
.A2(n_1311),
.B(n_1307),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1214),
.B(n_1281),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1281),
.A2(n_1198),
.B1(n_1202),
.B2(n_1200),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1247),
.B(n_1287),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1185),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1185),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1247),
.B(n_1287),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1247),
.B(n_1287),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1294),
.A2(n_1198),
.B(n_1200),
.C(n_1185),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1247),
.B(n_1287),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1217),
.A2(n_1198),
.B(n_1200),
.C(n_1185),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1296),
.A2(n_1198),
.B1(n_1202),
.B2(n_1200),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1216),
.A2(n_1198),
.B(n_1185),
.Y(n_1402)
);

O2A1O1Ixp5_ASAP7_75t_L g1403 ( 
.A1(n_1294),
.A2(n_1286),
.B(n_1319),
.C(n_1215),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1185),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1322),
.A2(n_1198),
.B(n_1185),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1231),
.A2(n_1242),
.B(n_1224),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1294),
.A2(n_1286),
.B(n_1319),
.C(n_1215),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1264),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1229),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1331),
.Y(n_1411)
);

INVxp67_ASAP7_75t_R g1412 ( 
.A(n_1380),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1387),
.B(n_1365),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1326),
.B(n_1408),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1348),
.A2(n_1400),
.B1(n_1359),
.B2(n_1360),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1365),
.B(n_1338),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1388),
.A2(n_1398),
.A3(n_1352),
.B(n_1404),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1379),
.A2(n_1353),
.B(n_1383),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1390),
.B(n_1396),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1399),
.B(n_1401),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1325),
.B(n_1332),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1365),
.B(n_1406),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1355),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1356),
.B(n_1389),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1365),
.B(n_1350),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1359),
.B(n_1393),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1330),
.A2(n_1343),
.B(n_1347),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1350),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1356),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1350),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1349),
.A2(n_1337),
.B(n_1357),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1343),
.B(n_1394),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1402),
.B(n_1384),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1398),
.A2(n_1405),
.B(n_1391),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1397),
.B(n_1328),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1327),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1358),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1382),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1376),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1328),
.B(n_1335),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1382),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1376),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1329),
.B(n_1363),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1329),
.B(n_1363),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1392),
.A2(n_1381),
.B(n_1339),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1403),
.B(n_1407),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1403),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1395),
.A2(n_1385),
.B(n_1340),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1341),
.B(n_1375),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1361),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1382),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1441),
.B(n_1372),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1452),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1433),
.B(n_1366),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1416),
.A2(n_1336),
.B1(n_1407),
.B2(n_1409),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1425),
.B(n_1386),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1435),
.A2(n_1370),
.B1(n_1373),
.B2(n_1354),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1411),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1417),
.B(n_1333),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1426),
.B(n_1334),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1440),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1423),
.B(n_1333),
.Y(n_1465)
);

NAND2x1_ASAP7_75t_L g1466 ( 
.A(n_1423),
.B(n_1378),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1345),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1435),
.A2(n_1346),
.B1(n_1351),
.B2(n_1368),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1429),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1431),
.A2(n_1330),
.B(n_1347),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1410),
.B(n_1342),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1424),
.Y(n_1473)
);

OAI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1432),
.A2(n_1434),
.B1(n_1447),
.B2(n_1444),
.C(n_1445),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1415),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1455),
.A2(n_1431),
.B(n_1419),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1467),
.B(n_1411),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1461),
.B(n_1369),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_R g1479 ( 
.A(n_1461),
.B(n_1364),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1467),
.B(n_1425),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1466),
.B(n_1414),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1454),
.A2(n_1449),
.B1(n_1435),
.B2(n_1446),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1466),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1454),
.A2(n_1449),
.B1(n_1435),
.B2(n_1446),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1410),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1473),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1466),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1464),
.Y(n_1489)
);

OA222x2_ASAP7_75t_L g1490 ( 
.A1(n_1474),
.A2(n_1434),
.B1(n_1414),
.B2(n_1450),
.C1(n_1441),
.C2(n_1448),
.Y(n_1490)
);

NAND4xp25_ASAP7_75t_L g1491 ( 
.A(n_1474),
.B(n_1447),
.C(n_1441),
.D(n_1444),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1465),
.A2(n_1449),
.B1(n_1446),
.B2(n_1445),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1465),
.A2(n_1447),
.B1(n_1444),
.B2(n_1445),
.C(n_1448),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1465),
.B(n_1414),
.Y(n_1494)
);

OAI211xp5_ASAP7_75t_L g1495 ( 
.A1(n_1457),
.A2(n_1436),
.B(n_1428),
.C(n_1450),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

NAND4xp25_ASAP7_75t_L g1498 ( 
.A(n_1457),
.B(n_1436),
.C(n_1450),
.D(n_1440),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1462),
.A2(n_1434),
.B1(n_1427),
.B2(n_1414),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1459),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1460),
.A2(n_1449),
.B1(n_1446),
.B2(n_1434),
.Y(n_1501)
);

AOI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1469),
.A2(n_1427),
.B1(n_1438),
.B2(n_1420),
.C1(n_1421),
.C2(n_1443),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1469),
.A2(n_1434),
.B1(n_1414),
.B2(n_1422),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1456),
.B(n_1451),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1475),
.B(n_1458),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_R g1506 ( 
.A(n_1472),
.B(n_1371),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1473),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1463),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1487),
.Y(n_1509)
);

INVx4_ASAP7_75t_SL g1510 ( 
.A(n_1481),
.Y(n_1510)
);

OR2x2_ASAP7_75t_SL g1511 ( 
.A(n_1490),
.B(n_1470),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1492),
.B(n_1413),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_SL g1513 ( 
.A(n_1495),
.B(n_1443),
.C(n_1460),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1493),
.A2(n_1439),
.B(n_1442),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_R g1516 ( 
.A(n_1478),
.B(n_1368),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1493),
.B(n_1463),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1476),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1497),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1497),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1476),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1476),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1505),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1497),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1481),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1482),
.A2(n_1442),
.B(n_1439),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1483),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1453),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1498),
.A2(n_1434),
.B(n_1418),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1453),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1483),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1525),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1515),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1523),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1523),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1486),
.Y(n_1539)
);

NAND4xp25_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1491),
.C(n_1495),
.D(n_1485),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1517),
.B(n_1531),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1512),
.B(n_1506),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.B(n_1488),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1509),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1513),
.A2(n_1498),
.B(n_1491),
.C(n_1489),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1509),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1489),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1533),
.B(n_1490),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1510),
.B(n_1532),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1514),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1486),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1534),
.B(n_1477),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1477),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1532),
.A2(n_1501),
.B1(n_1502),
.B2(n_1412),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1526),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1516),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1532),
.A2(n_1503),
.B(n_1499),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1525),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1515),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1534),
.B(n_1484),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1548),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1548),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1536),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1526),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1536),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1551),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1526),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1559),
.B(n_1510),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1540),
.A2(n_1515),
.B1(n_1525),
.B2(n_1519),
.C(n_1520),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1551),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1559),
.A2(n_1512),
.B1(n_1515),
.B2(n_1529),
.Y(n_1588)
);

OAI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1540),
.A2(n_1512),
.B(n_1502),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1553),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1564),
.B(n_1515),
.Y(n_1591)
);

AO21x1_ASAP7_75t_L g1592 ( 
.A1(n_1549),
.A2(n_1573),
.B(n_1542),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1512),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1571),
.B(n_1510),
.Y(n_1595)
);

XNOR2xp5_ASAP7_75t_L g1596 ( 
.A(n_1571),
.B(n_1511),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1544),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1564),
.B(n_1515),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1541),
.B(n_1504),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1545),
.B(n_1484),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1545),
.B(n_1534),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1569),
.A2(n_1575),
.B1(n_1536),
.B2(n_1561),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1563),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1504),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.B(n_1472),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

NAND2x1_ASAP7_75t_L g1611 ( 
.A(n_1565),
.B(n_1534),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1578),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1595),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1589),
.B(n_1535),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1609),
.B(n_1556),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1588),
.A2(n_1586),
.B1(n_1593),
.B2(n_1569),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1595),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1608),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1602),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1603),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1603),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1596),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1574),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1577),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1602),
.Y(n_1625)
);

AO22x1_ASAP7_75t_L g1626 ( 
.A1(n_1585),
.A2(n_1560),
.B1(n_1561),
.B2(n_1575),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1579),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1583),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1587),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1597),
.B(n_1558),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1581),
.B(n_1537),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1588),
.A2(n_1575),
.B1(n_1572),
.B2(n_1525),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1631),
.B(n_1558),
.Y(n_1637)
);

AOI21xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1616),
.A2(n_1544),
.B(n_1530),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1612),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1630),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1636),
.B(n_1606),
.C(n_1572),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1625),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1630),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1611),
.C(n_1591),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1636),
.A2(n_1585),
.B1(n_1560),
.B2(n_1598),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1620),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_R g1648 ( 
.A(n_1614),
.B(n_1560),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1623),
.A2(n_1582),
.B(n_1580),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1623),
.A2(n_1511),
.B1(n_1544),
.B2(n_1585),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1613),
.B(n_1599),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1566),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1617),
.A2(n_1582),
.B(n_1580),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1622),
.A2(n_1610),
.B1(n_1519),
.B2(n_1520),
.C(n_1525),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1619),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1639),
.B(n_1637),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1641),
.A2(n_1560),
.B1(n_1610),
.B2(n_1520),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1642),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_R g1661 ( 
.A(n_1653),
.B(n_1632),
.Y(n_1661)
);

INVx4_ASAP7_75t_L g1662 ( 
.A(n_1640),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1654),
.B(n_1618),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1648),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1652),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1650),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1662),
.B(n_1644),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_SL g1668 ( 
.A(n_1657),
.B(n_1638),
.C(n_1645),
.D(n_1655),
.Y(n_1668)
);

OAI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1660),
.A2(n_1643),
.B(n_1649),
.C(n_1646),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1663),
.A2(n_1511),
.B1(n_1628),
.B2(n_1615),
.Y(n_1670)
);

AO221x1_ASAP7_75t_L g1671 ( 
.A1(n_1664),
.A2(n_1651),
.B1(n_1634),
.B2(n_1647),
.C(n_1648),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1659),
.A2(n_1626),
.B(n_1633),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1520),
.B1(n_1519),
.B2(n_1529),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1658),
.A2(n_1635),
.B1(n_1629),
.B2(n_1627),
.C(n_1624),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1656),
.B(n_1632),
.C(n_1565),
.D(n_1607),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1666),
.B(n_1566),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1672),
.A2(n_1670),
.B1(n_1668),
.B2(n_1669),
.C(n_1674),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1667),
.B(n_1662),
.C(n_1520),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1671),
.A2(n_1605),
.B(n_1604),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1677),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1673),
.A2(n_1519),
.B1(n_1543),
.B2(n_1547),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_L g1683 ( 
.A(n_1678),
.B(n_1675),
.C(n_1676),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1681),
.B(n_1537),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1679),
.B(n_1538),
.C(n_1519),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1680),
.B(n_1538),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1682),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1681),
.B(n_1567),
.Y(n_1688)
);

NAND2xp33_ASAP7_75t_R g1689 ( 
.A(n_1686),
.B(n_1543),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1683),
.A2(n_1543),
.B1(n_1547),
.B2(n_1562),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1688),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1687),
.B(n_1528),
.C(n_1344),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1684),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1693),
.B(n_1685),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1691),
.B(n_1690),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1689),
.A2(n_1543),
.B1(n_1562),
.B2(n_1547),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1695),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1694),
.B1(n_1696),
.B2(n_1692),
.Y(n_1698)
);

OAI22x1_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1697),
.B1(n_1530),
.B2(n_1562),
.Y(n_1699)
);

OAI22x1_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1530),
.B1(n_1562),
.B2(n_1547),
.Y(n_1700)
);

AO22x2_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1563),
.B1(n_1530),
.B2(n_1568),
.Y(n_1701)
);

NAND3x1_ASAP7_75t_L g1702 ( 
.A(n_1701),
.B(n_1568),
.C(n_1576),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1527),
.B1(n_1522),
.B2(n_1518),
.Y(n_1703)
);

AO21x2_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1576),
.B(n_1567),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1552),
.B(n_1550),
.Y(n_1705)
);

AOI22x1_ASAP7_75t_L g1706 ( 
.A1(n_1704),
.A2(n_1546),
.B1(n_1550),
.B2(n_1552),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1705),
.A2(n_1518),
.B1(n_1522),
.B2(n_1527),
.C(n_1521),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1706),
.B(n_1546),
.C(n_1527),
.Y(n_1708)
);


endmodule