module fake_aes_5308_n_805 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_805);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_805;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_228;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_134;
wire n_656;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_19), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_78), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_85), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_45), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_26), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_18), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_102), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_103), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_89), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_47), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_91), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_57), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_39), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_74), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_41), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_28), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_80), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_36), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_53), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_10), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_40), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_42), .Y(n_134) );
CKINVDCx14_ASAP7_75t_R g135 ( .A(n_5), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_46), .B(n_93), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_58), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_73), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_20), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_48), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_44), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_70), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_25), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_8), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_129), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_121), .B(n_0), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_129), .B(n_0), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_131), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_152) );
OAI22x1_ASAP7_75t_SL g153 ( .A1(n_131), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_105), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_138), .B(n_4), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
INVx5_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_105), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_110), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_106), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_106), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_113), .A2(n_56), .B(n_101), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_116), .B(n_6), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_107), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_114), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_150), .B(n_115), .Y(n_171) );
AOI21x1_ASAP7_75t_L g172 ( .A1(n_164), .A2(n_139), .B(n_145), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_149), .B(n_117), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
AND3x2_ASAP7_75t_L g175 ( .A(n_150), .B(n_146), .C(n_122), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_154), .B(n_107), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_154), .B(n_119), .Y(n_180) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_155), .B(n_124), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_155), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_149), .B(n_126), .Y(n_188) );
AOI21x1_ASAP7_75t_L g189 ( .A1(n_164), .A2(n_144), .B(n_142), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_161), .B(n_111), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_158), .B(n_133), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_155), .Y(n_195) );
INVx8_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_166), .B(n_111), .Y(n_199) );
BUFx6f_ASAP7_75t_SL g200 ( .A(n_159), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_192), .B(n_161), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_192), .B(n_159), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_181), .A2(n_165), .B1(n_152), .B2(n_148), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_196), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_177), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_180), .B(n_159), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_171), .B(n_160), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_199), .B(n_160), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_181), .B(n_160), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_195), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_181), .A2(n_165), .B1(n_148), .B2(n_156), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_195), .B(n_162), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_194), .B(n_162), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_195), .B(n_162), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_195), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_197), .B(n_165), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVxp67_ASAP7_75t_SL g219 ( .A(n_187), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_187), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_187), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_197), .B(n_112), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_196), .B(n_112), .Y(n_223) );
NAND3xp33_ASAP7_75t_L g224 ( .A(n_185), .B(n_156), .C(n_152), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_196), .A2(n_132), .B1(n_156), .B2(n_130), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_183), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_173), .B(n_130), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_168), .B(n_137), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_168), .Y(n_230) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_173), .B(n_134), .C(n_141), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_168), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_188), .B(n_137), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_169), .A2(n_153), .B1(n_140), .B2(n_143), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_188), .B(n_140), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_196), .B(n_143), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_196), .B(n_118), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_200), .B(n_120), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_169), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_184), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_169), .B(n_123), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_191), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g245 ( .A(n_185), .B(n_125), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_191), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g247 ( .A(n_185), .B(n_127), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_169), .B(n_128), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_186), .B(n_193), .C(n_201), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_218), .A2(n_193), .B(n_186), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_227), .B(n_175), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_226), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_227), .B(n_233), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_239), .B(n_200), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_239), .B(n_200), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_208), .B(n_175), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_218), .A2(n_193), .B(n_186), .Y(n_257) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_204), .A2(n_193), .B(n_186), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_206), .B(n_153), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_164), .B(n_198), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_233), .B(n_114), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_232), .A2(n_172), .B(n_189), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_240), .A2(n_198), .B(n_201), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_240), .A2(n_172), .B(n_189), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_217), .A2(n_136), .B(n_167), .C(n_114), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_207), .A2(n_200), .B(n_198), .C(n_190), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_235), .B(n_7), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_204), .A2(n_167), .B1(n_157), .B2(n_179), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_235), .B(n_167), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_243), .A2(n_190), .B(n_170), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_241), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_241), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_230), .A2(n_190), .B(n_170), .Y(n_276) );
AO21x1_ASAP7_75t_L g277 ( .A1(n_231), .A2(n_170), .B(n_174), .Y(n_277) );
AO21x1_ASAP7_75t_L g278 ( .A1(n_229), .A2(n_174), .B(n_176), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_248), .A2(n_179), .B(n_178), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_241), .B(n_157), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_210), .B(n_7), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_228), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_209), .B(n_8), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_205), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_203), .A2(n_167), .B(n_157), .C(n_178), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_211), .A2(n_179), .B(n_178), .Y(n_286) );
AOI21x1_ASAP7_75t_L g287 ( .A1(n_223), .A2(n_176), .B(n_174), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_250), .A2(n_216), .B(n_211), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_257), .A2(n_247), .B(n_245), .Y(n_289) );
AOI21x1_ASAP7_75t_L g290 ( .A1(n_260), .A2(n_246), .B(n_244), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_265), .A2(n_213), .B(n_215), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_270), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_265), .A2(n_246), .B(n_244), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_263), .A2(n_236), .B(n_222), .Y(n_294) );
OAI22x1_ASAP7_75t_L g295 ( .A1(n_259), .A2(n_234), .B1(n_224), .B2(n_214), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_264), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_262), .A2(n_246), .B(n_244), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_258), .A2(n_224), .B(n_237), .C(n_228), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_273), .A2(n_216), .B(n_219), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g300 ( .A1(n_252), .A2(n_242), .B(n_237), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_276), .A2(n_216), .B(n_221), .Y(n_301) );
CKINVDCx6p67_ASAP7_75t_R g302 ( .A(n_274), .Y(n_302) );
OAI21x1_ASAP7_75t_SL g303 ( .A1(n_267), .A2(n_242), .B(n_237), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_278), .A2(n_242), .B(n_228), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_253), .B(n_212), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_274), .B(n_205), .Y(n_306) );
AOI221xp5_ASAP7_75t_SL g307 ( .A1(n_249), .A2(n_225), .B1(n_221), .B2(n_220), .C(n_238), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_251), .B(n_234), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_221), .B(n_220), .C(n_157), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_275), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_274), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_256), .B(n_220), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_274), .B(n_9), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_302), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_303), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_305), .B(n_271), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_287), .B(n_254), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_293), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_297), .A2(n_255), .B(n_277), .Y(n_321) );
OR3x4_ASAP7_75t_SL g322 ( .A(n_295), .B(n_10), .C(n_11), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_310), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_308), .B(n_283), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_296), .B(n_269), .Y(n_326) );
AO31x2_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_266), .A3(n_285), .B(n_261), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_290), .A2(n_279), .B(n_276), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_302), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_298), .B(n_281), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_291), .A2(n_268), .B(n_272), .Y(n_332) );
NOR2xp33_ASAP7_75t_R g333 ( .A(n_311), .B(n_275), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_294), .A2(n_286), .B(n_280), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_307), .A2(n_309), .B(n_301), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_315), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
AO21x1_ASAP7_75t_SL g340 ( .A1(n_320), .A2(n_313), .B(n_312), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_317), .A2(n_292), .B1(n_309), .B2(n_306), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_326), .B(n_306), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_314), .B(n_275), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_289), .B(n_299), .Y(n_349) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_316), .B(n_284), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_333), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_284), .B1(n_157), .B2(n_176), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_334), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_324), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_317), .B(n_284), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_331), .B(n_11), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_329), .B(n_12), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_326), .B(n_12), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_356), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_338), .B(n_321), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_338), .B(n_336), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_342), .B(n_336), .Y(n_379) );
AO31x2_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_330), .A3(n_335), .B(n_331), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_352), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_361), .B(n_329), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_342), .B(n_336), .Y(n_384) );
OR2x6_ASAP7_75t_L g385 ( .A(n_345), .B(n_321), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_361), .B(n_337), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_370), .B(n_335), .C(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_352), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_372), .B(n_336), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_359), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_343), .B(n_336), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_321), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_372), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_357), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_344), .B(n_327), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_347), .B(n_319), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_347), .B(n_327), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_327), .Y(n_404) );
INVx4_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_327), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_364), .B(n_327), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_364), .B(n_327), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_355), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_332), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_339), .B(n_332), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_368), .A2(n_332), .B1(n_322), .B2(n_157), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_363), .B(n_332), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_369), .B(n_13), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_157), .B1(n_182), .B2(n_15), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_13), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_366), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_339), .B(n_14), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_339), .B(n_15), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_341), .B(n_16), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_341), .B(n_16), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_341), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_404), .B(n_366), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_373), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_419), .B(n_353), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_376), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_419), .B(n_353), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_376), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_396), .A2(n_366), .B1(n_362), .B2(n_341), .C1(n_353), .C2(n_358), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_377), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_404), .B(n_362), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_421), .B(n_362), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_402), .B(n_353), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_373), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_377), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_400), .B(n_362), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_400), .B(n_371), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_383), .B(n_349), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_399), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_403), .B(n_411), .Y(n_449) );
OAI22xp33_ASAP7_75t_SL g450 ( .A1(n_387), .A2(n_348), .B1(n_350), .B2(n_367), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_387), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_387), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_419), .B(n_371), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_381), .Y(n_455) );
NAND2x1p5_ASAP7_75t_SL g456 ( .A(n_415), .B(n_350), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_419), .B(n_393), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_420), .A2(n_340), .B1(n_349), .B2(n_371), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_403), .B(n_367), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_383), .B(n_349), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_381), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_411), .B(n_367), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_382), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_382), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_389), .A2(n_340), .B1(n_349), .B2(n_348), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_390), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_412), .B(n_348), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_412), .B(n_17), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_390), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_386), .B(n_17), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_386), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_413), .B(n_21), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_422), .A2(n_22), .B(n_23), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_388), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_405), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_393), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_397), .B(n_24), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_373), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_375), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_426), .B(n_27), .C(n_29), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_375), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_413), .B(n_30), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_397), .B(n_31), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_405), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_378), .B(n_32), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_378), .B(n_34), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_379), .B(n_384), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_375), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_398), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_424), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_408), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_379), .B(n_35), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_385), .A2(n_182), .B1(n_38), .B2(n_43), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_408), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_384), .B(n_37), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_392), .B(n_49), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_398), .B(n_50), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_406), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_394), .B(n_51), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_394), .B(n_52), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_385), .A2(n_182), .B1(n_55), .B2(n_59), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_418), .B(n_54), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_374), .B(n_60), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_410), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_424), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_410), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_406), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_418), .B(n_61), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_385), .A2(n_429), .B1(n_423), .B2(n_430), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_407), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_407), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_374), .B(n_63), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_380), .B(n_64), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_395), .B(n_65), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_429), .B(n_66), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_395), .B(n_68), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_414), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_449), .B(n_409), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_435), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_449), .B(n_409), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_435), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_437), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_517), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_437), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_487), .B(n_409), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_487), .B(n_415), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_461), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_471), .B(n_380), .Y(n_528) );
BUFx2_ASAP7_75t_SL g529 ( .A(n_451), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_468), .B(n_380), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_467), .B(n_405), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_440), .B(n_385), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_478), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_461), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_440), .B(n_385), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_468), .B(n_380), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_490), .B(n_380), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_448), .B(n_380), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_445), .B(n_374), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_445), .B(n_374), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_432), .B(n_401), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_479), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_475), .Y(n_543) );
AND3x2_ASAP7_75t_L g544 ( .A(n_433), .B(n_401), .C(n_428), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_488), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_467), .B(n_405), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_463), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_455), .B(n_416), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_463), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_476), .B(n_416), .Y(n_550) );
AND2x4_ASAP7_75t_SL g551 ( .A(n_451), .B(n_431), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_464), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_464), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_433), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_466), .Y(n_555) );
INVxp67_ASAP7_75t_R g556 ( .A(n_514), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_466), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_469), .B(n_425), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_469), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_489), .B(n_425), .Y(n_560) );
NAND2x1_ASAP7_75t_L g561 ( .A(n_475), .B(n_431), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_457), .B(n_401), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_432), .B(n_401), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_443), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_498), .Y(n_566) );
AND2x4_ASAP7_75t_SL g567 ( .A(n_475), .B(n_427), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_498), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_505), .B(n_427), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_457), .B(n_427), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_517), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_452), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_439), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_446), .B(n_417), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_511), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_442), .B(n_417), .Y(n_576) );
BUFx2_ASAP7_75t_L g577 ( .A(n_484), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_452), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_457), .B(n_427), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_481), .B(n_414), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_470), .A2(n_391), .B1(n_182), .B2(n_72), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_511), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_507), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_439), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_446), .B(n_391), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_510), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_447), .B(n_391), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_459), .B(n_391), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_444), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_444), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_484), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_459), .B(n_391), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_484), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_438), .B(n_182), .C(n_71), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_462), .B(n_69), .Y(n_595) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_513), .B(n_75), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_462), .B(n_77), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_454), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_434), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_509), .A2(n_182), .B1(n_81), .B2(n_82), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_460), .B(n_79), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_502), .B(n_83), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_454), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_474), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_474), .Y(n_605) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_450), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_502), .B(n_86), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_441), .B(n_87), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_491), .Y(n_609) );
NOR2x1p5_ASAP7_75t_SL g610 ( .A(n_513), .B(n_88), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_508), .B(n_90), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_434), .B(n_92), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g613 ( .A(n_561), .B(n_508), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_563), .B(n_543), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_525), .B(n_436), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_574), .B(n_441), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_526), .B(n_491), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_528), .B(n_504), .Y(n_618) );
NAND2xp33_ASAP7_75t_SL g619 ( .A(n_577), .B(n_512), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_518), .B(n_504), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
AND2x2_ASAP7_75t_SL g622 ( .A(n_596), .B(n_512), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_538), .B(n_506), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_529), .B(n_512), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_571), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_596), .A2(n_465), .B(n_503), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_530), .B(n_482), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_586), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_533), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_536), .B(n_482), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_520), .B(n_436), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_539), .B(n_436), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_533), .Y(n_634) );
NAND2x1_ASAP7_75t_L g635 ( .A(n_543), .B(n_503), .Y(n_635) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_554), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_545), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_606), .A2(n_458), .B(n_501), .C(n_493), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_606), .B(n_494), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_545), .B(n_472), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_576), .B(n_494), .Y(n_641) );
OAI21xp33_ASAP7_75t_SL g642 ( .A1(n_543), .A2(n_516), .B(n_514), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_591), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_563), .B(n_434), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_542), .B(n_506), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_580), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_521), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_522), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_524), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_527), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_534), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_547), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_566), .B(n_453), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_573), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_594), .B(n_480), .C(n_516), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_568), .B(n_453), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_572), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_573), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_539), .B(n_453), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_542), .B(n_472), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_549), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_572), .B(n_456), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_540), .B(n_503), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_552), .B(n_495), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_578), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_612), .B(n_495), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_553), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_555), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_575), .B(n_492), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_540), .B(n_500), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_601), .B(n_473), .C(n_515), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_563), .B(n_500), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_599), .B(n_486), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_541), .B(n_499), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g677 ( .A(n_565), .B(n_477), .C(n_483), .D(n_497), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_582), .B(n_499), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_557), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_559), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_554), .Y(n_681) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_565), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_541), .B(n_492), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_532), .A2(n_486), .B1(n_485), .B2(n_496), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_564), .B(n_485), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_584), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_562), .B(n_456), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_578), .B(n_496), .Y(n_688) );
NOR2x1p5_ASAP7_75t_L g689 ( .A(n_537), .B(n_94), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_569), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_616), .B(n_599), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_639), .B(n_523), .Y(n_692) );
OAI222xp33_ASAP7_75t_L g693 ( .A1(n_624), .A2(n_531), .B1(n_546), .B2(n_535), .C1(n_532), .C2(n_570), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_626), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_690), .B(n_551), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_642), .A2(n_556), .B1(n_535), .B2(n_579), .Y(n_696) );
NOR2x1_ASAP7_75t_R g697 ( .A(n_682), .B(n_612), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_661), .B(n_585), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_634), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_615), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_629), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_645), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_649), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_642), .A2(n_588), .B1(n_592), .B2(n_600), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_622), .A2(n_600), .B1(n_551), .B2(n_607), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_681), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_639), .B(n_523), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_646), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_650), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_651), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_652), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_653), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_620), .B(n_587), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_618), .B(n_604), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_641), .B(n_589), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_668), .A2(n_567), .B1(n_612), .B2(n_597), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_617), .B(n_598), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_618), .B(n_605), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_623), .B(n_590), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_633), .B(n_567), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_621), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_625), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_654), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_663), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_669), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_632), .B(n_544), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_670), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_623), .B(n_603), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_679), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_644), .B(n_544), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_613), .A2(n_610), .B(n_611), .C(n_602), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_680), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_624), .Y(n_733) );
OAI32xp33_ASAP7_75t_L g734 ( .A1(n_619), .A2(n_595), .A3(n_608), .B1(n_550), .B2(n_548), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_655), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_655), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_630), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_637), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_695), .B(n_667), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_696), .A2(n_638), .B1(n_624), .B2(n_657), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_708), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_733), .A2(n_627), .B(n_635), .C(n_657), .Y(n_742) );
OA22x2_ASAP7_75t_L g743 ( .A1(n_733), .A2(n_614), .B1(n_644), .B2(n_674), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_692), .B(n_648), .Y(n_744) );
OAI21xp33_ASAP7_75t_L g745 ( .A1(n_704), .A2(n_664), .B(n_636), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_705), .A2(n_668), .B1(n_716), .B2(n_700), .Y(n_746) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_730), .Y(n_747) );
OAI31xp33_ASAP7_75t_L g748 ( .A1(n_693), .A2(n_689), .A3(n_614), .B(n_659), .Y(n_748) );
AOI31xp33_ASAP7_75t_L g749 ( .A1(n_697), .A2(n_684), .A3(n_688), .B(n_674), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_734), .A2(n_677), .B1(n_687), .B2(n_658), .C(n_631), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_716), .A2(n_675), .B1(n_662), .B2(n_673), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_714), .Y(n_752) );
NOR2xp67_ASAP7_75t_L g753 ( .A(n_726), .B(n_647), .Y(n_753) );
AOI21xp33_ASAP7_75t_SL g754 ( .A1(n_731), .A2(n_677), .B(n_643), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_699), .A2(n_675), .B1(n_640), .B2(n_628), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_708), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_692), .A2(n_687), .B(n_658), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_735), .A2(n_665), .B1(n_672), .B2(n_683), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_714), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g760 ( .A1(n_720), .A2(n_676), .B(n_685), .C(n_678), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_694), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_706), .A2(n_581), .B(n_678), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_707), .B(n_581), .C(n_608), .Y(n_763) );
AO21x1_ASAP7_75t_L g764 ( .A1(n_701), .A2(n_671), .B(n_666), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_747), .B(n_736), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_754), .A2(n_707), .B1(n_732), .B2(n_729), .C(n_703), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_754), .A2(n_709), .B1(n_702), .B2(n_727), .C(n_725), .Y(n_767) );
AOI211xp5_ASAP7_75t_L g768 ( .A1(n_746), .A2(n_710), .B(n_711), .C(n_724), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_744), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_749), .A2(n_712), .B1(n_723), .B2(n_718), .C(n_728), .Y(n_770) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_745), .A2(n_718), .B1(n_728), .B2(n_737), .C(n_738), .Y(n_771) );
AOI21xp33_ASAP7_75t_L g772 ( .A1(n_748), .A2(n_719), .B(n_671), .Y(n_772) );
NAND2x1_ASAP7_75t_L g773 ( .A(n_753), .B(n_698), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_740), .A2(n_691), .B(n_721), .C(n_722), .Y(n_774) );
INVxp67_ASAP7_75t_SL g775 ( .A(n_741), .Y(n_775) );
AO22x1_ASAP7_75t_L g776 ( .A1(n_756), .A2(n_686), .B1(n_660), .B2(n_656), .Y(n_776) );
NAND4xp25_ASAP7_75t_L g777 ( .A(n_742), .B(n_750), .C(n_751), .D(n_739), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_743), .A2(n_715), .B(n_717), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_769), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_770), .B(n_764), .Y(n_780) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_777), .B(n_763), .C(n_762), .D(n_757), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_774), .B(n_761), .C(n_755), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g783 ( .A1(n_768), .A2(n_759), .B(n_752), .Y(n_783) );
NOR2x1_ASAP7_75t_L g784 ( .A(n_773), .B(n_760), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_765), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_785), .B(n_775), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_781), .B(n_772), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_784), .B(n_778), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_782), .B(n_771), .Y(n_789) );
NOR2x1p5_ASAP7_75t_L g790 ( .A(n_786), .B(n_779), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g791 ( .A(n_789), .B(n_780), .C(n_767), .D(n_766), .Y(n_791) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_788), .B(n_783), .C(n_758), .D(n_776), .Y(n_792) );
NOR2x1_ASAP7_75t_L g793 ( .A(n_792), .B(n_787), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_790), .A2(n_713), .B(n_609), .C(n_584), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_794), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_793), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_796), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_795), .A2(n_791), .B1(n_560), .B2(n_558), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_797), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_799), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_800), .A2(n_798), .B(n_96), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_801), .Y(n_802) );
OA21x2_ASAP7_75t_L g803 ( .A1(n_802), .A2(n_95), .B(n_97), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_803), .B(n_98), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_804), .A2(n_99), .B1(n_100), .B2(n_104), .Y(n_805) );
endmodule