module fake_jpeg_11067_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_25),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_73),
.Y(n_93)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_99),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_70),
.B1(n_61),
.B2(n_64),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_84),
.B(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_66),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_72),
.B(n_58),
.C(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_50),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_69),
.C(n_77),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_6),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_88),
.B1(n_89),
.B2(n_61),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_65),
.B1(n_62),
.B2(n_52),
.Y(n_133)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_114),
.Y(n_152)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_127),
.B1(n_113),
.B2(n_108),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_55),
.B1(n_75),
.B2(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_127),
.B1(n_23),
.B2(n_46),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_73),
.B1(n_53),
.B2(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_135),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_64),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_133),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_7),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_2),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_149),
.B(n_9),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_53),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_3),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_4),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_8),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_6),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_131),
.CI(n_144),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_141),
.B1(n_150),
.B2(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_169),
.B1(n_10),
.B2(n_11),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx6p67_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_148),
.B1(n_11),
.B2(n_10),
.C(n_13),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_186),
.B1(n_175),
.B2(n_173),
.Y(n_188)
);

OAI322xp33_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_162),
.A3(n_153),
.B1(n_170),
.B2(n_157),
.C1(n_20),
.C2(n_22),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_175),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_190),
.A2(n_187),
.B(n_174),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_180),
.B1(n_182),
.B2(n_172),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_189),
.B(n_28),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_189),
.C(n_29),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_18),
.B(n_30),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_32),
.Y(n_197)
);


endmodule