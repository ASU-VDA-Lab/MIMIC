module fake_jpeg_3203_n_723 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_723);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_723;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_722;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_721;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_133),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_70),
.Y(n_203)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_71),
.Y(n_164)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_29),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_46),
.B(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_91),
.B(n_92),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_97),
.B(n_100),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_29),
.B(n_16),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_33),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_104),
.B(n_105),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_43),
.B(n_16),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_49),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_126),
.B(n_55),
.Y(n_181)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_38),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_56),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_32),
.B(n_15),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_35),
.B(n_58),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_136),
.B(n_140),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_71),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_142),
.B(n_181),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_49),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_150),
.B(n_155),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_51),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_152),
.B(n_221),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_55),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_60),
.B1(n_37),
.B2(n_41),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_163),
.A2(n_194),
.B1(n_200),
.B2(n_212),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_125),
.A2(n_56),
.B1(n_51),
.B2(n_44),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_179),
.A2(n_188),
.B1(n_209),
.B2(n_113),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_106),
.B(n_50),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_50),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_108),
.A2(n_56),
.B1(n_47),
.B2(n_60),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_84),
.A2(n_60),
.B1(n_41),
.B2(n_48),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_199),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_78),
.A2(n_41),
.B1(n_48),
.B2(n_52),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_48),
.B1(n_52),
.B2(n_58),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_206),
.A2(n_226),
.B1(n_1),
.B2(n_2),
.Y(n_307)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_113),
.B(n_22),
.CON(n_208),
.SN(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_208),
.A2(n_22),
.B(n_1),
.C(n_2),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_120),
.A2(n_47),
.B1(n_39),
.B2(n_35),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_93),
.A2(n_39),
.B1(n_32),
.B2(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_72),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_225),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_107),
.B(n_15),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_61),
.A2(n_22),
.B1(n_14),
.B2(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_67),
.B(n_14),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_121),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_232),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g363 ( 
.A(n_233),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_149),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_234),
.Y(n_373)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_237),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_238),
.B(n_268),
.Y(n_362)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_246),
.Y(n_320)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_241),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_247),
.B(n_284),
.Y(n_321)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_248),
.Y(n_340)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_249),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_208),
.A2(n_121),
.B(n_120),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_250),
.B(n_279),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_166),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_256),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_166),
.A2(n_89),
.B1(n_96),
.B2(n_117),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_254),
.A2(n_273),
.B1(n_297),
.B2(n_299),
.Y(n_319)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_143),
.Y(n_255)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_166),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_191),
.A2(n_200),
.B1(n_135),
.B2(n_154),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_257),
.A2(n_280),
.B1(n_304),
.B2(n_307),
.Y(n_370)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_259),
.Y(n_361)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_137),
.Y(n_264)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVx6_ASAP7_75t_SL g338 ( 
.A(n_265),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_62),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_145),
.B(n_63),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_270),
.B(n_272),
.Y(n_375)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_141),
.B(n_10),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_205),
.A2(n_128),
.B1(n_123),
.B2(n_94),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx6_ASAP7_75t_SL g369 ( 
.A(n_274),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_176),
.Y(n_276)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_157),
.B(n_13),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_277),
.B(n_296),
.Y(n_330)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_212),
.A2(n_188),
.B1(n_65),
.B2(n_69),
.Y(n_280)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_283),
.Y(n_329)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_195),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_287),
.Y(n_332)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_147),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_170),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_289),
.Y(n_365)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_290),
.Y(n_313)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_291),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_179),
.A2(n_77),
.B1(n_74),
.B2(n_13),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_292),
.A2(n_298),
.B1(n_3),
.B2(n_5),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_152),
.B(n_174),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_293),
.B(n_295),
.Y(n_371)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_294),
.Y(n_357)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_164),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_158),
.B(n_12),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_168),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_160),
.B(n_12),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_164),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_151),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_229),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_162),
.Y(n_305)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_161),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_203),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_206),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_310),
.B1(n_221),
.B2(n_220),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_209),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_144),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_227),
.B1(n_218),
.B2(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_172),
.B(n_11),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_1),
.Y(n_334)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_323),
.A2(n_337),
.B1(n_348),
.B2(n_360),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_252),
.A2(n_138),
.B1(n_177),
.B2(n_192),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_326),
.A2(n_343),
.B1(n_344),
.B2(n_367),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_334),
.B(n_351),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_186),
.B1(n_220),
.B2(n_171),
.Y(n_337)
);

NAND2x2_ASAP7_75t_SL g339 ( 
.A(n_265),
.B(n_218),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g427 ( 
.A1(n_339),
.A2(n_7),
.B(n_8),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_250),
.A2(n_260),
.B1(n_308),
.B2(n_266),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_260),
.A2(n_161),
.B1(n_173),
.B2(n_182),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_230),
.A2(n_162),
.B1(n_186),
.B2(n_171),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_263),
.B(n_180),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_293),
.A2(n_227),
.B1(n_165),
.B2(n_215),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_267),
.A2(n_211),
.B1(n_223),
.B2(n_218),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_353),
.A2(n_368),
.B1(n_304),
.B2(n_269),
.Y(n_385)
);

AOI22x1_ASAP7_75t_L g355 ( 
.A1(n_267),
.A2(n_134),
.B1(n_190),
.B2(n_148),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_355),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_148),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_366),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_273),
.A2(n_182),
.B1(n_173),
.B2(n_134),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_235),
.B(n_203),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_281),
.A2(n_190),
.B1(n_5),
.B2(n_6),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_301),
.A2(n_190),
.B1(n_6),
.B2(n_7),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_288),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_251),
.B(n_3),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_7),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_370),
.A2(n_254),
.B1(n_305),
.B2(n_306),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_377),
.A2(n_381),
.B1(n_386),
.B2(n_392),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_244),
.C(n_231),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_384),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_382),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_370),
.A2(n_291),
.B1(n_262),
.B2(n_261),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_321),
.B(n_311),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_236),
.C(n_309),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_385),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_324),
.A2(n_264),
.B1(n_302),
.B2(n_233),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_387),
.B(n_388),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_303),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_389),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_369),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_402),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_324),
.A2(n_338),
.B1(n_327),
.B2(n_339),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_338),
.A2(n_300),
.B1(n_295),
.B2(n_237),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_333),
.B1(n_317),
.B2(n_358),
.Y(n_458)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_275),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_355),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_330),
.B(n_297),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_399),
.Y(n_449)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_289),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_327),
.A2(n_282),
.B1(n_299),
.B2(n_242),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_400),
.A2(n_360),
.B1(n_350),
.B2(n_313),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_339),
.A2(n_294),
.B1(n_290),
.B2(n_258),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_401),
.A2(n_405),
.B(n_416),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_274),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_239),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_403),
.B(n_404),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_249),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_327),
.A2(n_339),
.B(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_241),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_410),
.Y(n_447)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_415),
.B(n_418),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_345),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_419),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_345),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_421),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_424),
.Y(n_466)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_348),
.B(n_232),
.CI(n_259),
.CON(n_426),
.SN(n_426)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_380),
.A3(n_388),
.B1(n_397),
.B2(n_406),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_427),
.A2(n_9),
.B(n_376),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_392),
.A2(n_323),
.B(n_337),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_452),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_430),
.B(n_383),
.Y(n_482)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_355),
.B(n_367),
.C(n_319),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_437),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_414),
.A2(n_357),
.B1(n_313),
.B2(n_342),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_438),
.A2(n_458),
.B1(n_468),
.B2(n_422),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_417),
.A2(n_315),
.B1(n_372),
.B2(n_342),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_440),
.A2(n_441),
.B1(n_455),
.B2(n_381),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_417),
.A2(n_328),
.B1(n_357),
.B2(n_322),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_365),
.B(n_356),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_445),
.A2(n_448),
.B(n_450),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_401),
.A2(n_336),
.B(n_356),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_423),
.A2(n_336),
.B(n_314),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_376),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_424),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_391),
.A2(n_322),
.B1(n_347),
.B2(n_346),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_314),
.B(n_361),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_391),
.B(n_346),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_459),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_380),
.A2(n_347),
.B(n_333),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_462),
.B(n_398),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_335),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_384),
.C(n_415),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_394),
.B(n_317),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_467),
.B(n_410),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_377),
.A2(n_358),
.B1(n_335),
.B2(n_349),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

OAI32xp33_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_383),
.A3(n_403),
.B1(n_404),
.B2(n_399),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_472),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_451),
.A2(n_414),
.B1(n_425),
.B2(n_421),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_474),
.A2(n_489),
.B(n_446),
.Y(n_523)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_476),
.Y(n_522)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_477),
.Y(n_526)
);

XNOR2x1_ASAP7_75t_SL g478 ( 
.A(n_463),
.B(n_378),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_L g542 ( 
.A(n_478),
.B(n_482),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_393),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_479),
.Y(n_546)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_480),
.Y(n_528)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_483),
.A2(n_486),
.B(n_491),
.Y(n_530)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_484),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_465),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_373),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_487),
.A2(n_488),
.B1(n_493),
.B2(n_496),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_443),
.A2(n_426),
.B1(n_413),
.B2(n_387),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_490),
.A2(n_503),
.B1(n_440),
.B2(n_428),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_433),
.B(n_373),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_444),
.Y(n_492)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_492),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_428),
.A2(n_386),
.B1(n_426),
.B2(n_407),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_SL g494 ( 
.A(n_463),
.B(n_408),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_507),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_442),
.B(n_431),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_434),
.B(n_466),
.C(n_430),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_434),
.C(n_460),
.Y(n_511)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_469),
.Y(n_498)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_498),
.Y(n_549)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_500),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_409),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_502),
.Y(n_517)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_443),
.A2(n_395),
.B1(n_389),
.B2(n_419),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_467),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_506),
.Y(n_529)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_325),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_325),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_459),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_511),
.B(n_524),
.C(n_525),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_510),
.A2(n_451),
.B1(n_449),
.B2(n_464),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_513),
.A2(n_516),
.B1(n_534),
.B2(n_481),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_501),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_515),
.B(n_532),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_510),
.A2(n_451),
.B1(n_449),
.B2(n_464),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_504),
.A2(n_446),
.B(n_448),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_520),
.A2(n_523),
.B(n_535),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_521),
.A2(n_474),
.B1(n_481),
.B2(n_473),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_466),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_430),
.C(n_459),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_533),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_500),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_509),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_475),
.A2(n_429),
.B1(n_438),
.B2(n_468),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_504),
.A2(n_461),
.B(n_445),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g536 ( 
.A(n_506),
.B(n_436),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_536),
.B(n_450),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_490),
.A2(n_428),
.B1(n_441),
.B2(n_450),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_537),
.A2(n_493),
.B1(n_488),
.B2(n_495),
.Y(n_557)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_478),
.C(n_482),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_540),
.B(n_545),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_494),
.B(n_465),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_541),
.B(n_462),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_479),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_508),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_477),
.B(n_431),
.Y(n_544)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_544),
.Y(n_573)
);

XOR2x2_ASAP7_75t_L g545 ( 
.A(n_472),
.B(n_445),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_442),
.C(n_452),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_547),
.B(n_483),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_546),
.A2(n_475),
.B(n_495),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_551),
.A2(n_564),
.B(n_580),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_480),
.Y(n_552)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_552),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_505),
.Y(n_553)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_499),
.Y(n_555)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_517),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_566),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_557),
.A2(n_575),
.B1(n_582),
.B2(n_518),
.Y(n_602)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_558),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_561),
.A2(n_569),
.B1(n_576),
.B2(n_581),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

BUFx12f_ASAP7_75t_SL g564 ( 
.A(n_530),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_528),
.B(n_452),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_519),
.B(n_528),
.Y(n_568)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_544),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_513),
.B(n_476),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_570),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_529),
.B(n_471),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_577),
.Y(n_614)
);

A2O1A1Ixp33_ASAP7_75t_SL g607 ( 
.A1(n_572),
.A2(n_578),
.B(n_579),
.C(n_469),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g610 ( 
.A(n_574),
.B(n_340),
.C(n_349),
.Y(n_610)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_517),
.B(n_492),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_534),
.B(n_473),
.Y(n_578)
);

AO22x1_ASAP7_75t_SL g579 ( 
.A1(n_516),
.A2(n_503),
.B1(n_484),
.B2(n_437),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_523),
.A2(n_456),
.B(n_437),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_547),
.B(n_439),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_521),
.A2(n_456),
.B1(n_470),
.B2(n_458),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_520),
.A2(n_470),
.B(n_498),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_584),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_515),
.B(n_502),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_585),
.B(n_549),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_561),
.A2(n_519),
.B1(n_537),
.B2(n_514),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_586),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_570),
.A2(n_514),
.B1(n_535),
.B2(n_536),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_568),
.A2(n_536),
.B1(n_531),
.B2(n_539),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_550),
.A2(n_545),
.B1(n_541),
.B2(n_522),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_552),
.A2(n_512),
.B1(n_522),
.B2(n_538),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_594),
.B(n_613),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_550),
.A2(n_512),
.B1(n_548),
.B2(n_538),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_601),
.B1(n_603),
.B2(n_604),
.Y(n_638)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_598),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_573),
.A2(n_548),
.B1(n_542),
.B2(n_525),
.Y(n_601)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_602),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_573),
.A2(n_542),
.B1(n_527),
.B2(n_518),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_576),
.A2(n_439),
.B1(n_540),
.B2(n_511),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_557),
.A2(n_524),
.B1(n_432),
.B2(n_435),
.Y(n_605)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_605),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_432),
.C(n_361),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_606),
.B(n_611),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_607),
.A2(n_580),
.B(n_584),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_SL g619 ( 
.A(n_610),
.B(n_572),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_567),
.B(n_432),
.C(n_316),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_575),
.A2(n_419),
.B1(n_389),
.B2(n_411),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_612),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_616),
.B(n_618),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_608),
.A2(n_551),
.B(n_578),
.Y(n_617)
);

XNOR2x1_ASAP7_75t_L g660 ( 
.A(n_617),
.B(n_619),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_595),
.Y(n_618)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_592),
.Y(n_621)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_621),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_560),
.C(n_583),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_628),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_559),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_606),
.B(n_563),
.C(n_578),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_629),
.B(n_632),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_596),
.B(n_581),
.Y(n_630)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_630),
.Y(n_645)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_588),
.Y(n_631)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_631),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_605),
.B(n_563),
.C(n_571),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_601),
.B(n_602),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_633),
.B(n_590),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_566),
.Y(n_634)
);

OAI321xp33_ASAP7_75t_L g655 ( 
.A1(n_634),
.A2(n_553),
.A3(n_555),
.B1(n_565),
.B2(n_577),
.C(n_564),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_597),
.A2(n_554),
.B(n_572),
.Y(n_635)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_588),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_636),
.A2(n_558),
.B1(n_587),
.B2(n_556),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_637),
.B(n_615),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_596),
.B(n_574),
.C(n_579),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_639),
.B(n_640),
.C(n_600),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_608),
.B(n_579),
.C(n_565),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_612),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_641),
.A2(n_599),
.B1(n_589),
.B2(n_597),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_642),
.B(n_643),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_603),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_646),
.B(n_648),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_620),
.B(n_586),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_647),
.B(n_649),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_624),
.B(n_593),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_627),
.B(n_615),
.C(n_591),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_650),
.B(n_662),
.C(n_663),
.Y(n_673)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_652),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_653),
.A2(n_625),
.B1(n_631),
.B2(n_636),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_655),
.A2(n_607),
.B(n_585),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_579),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_659),
.B(n_661),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_638),
.B(n_614),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_622),
.B(n_582),
.C(n_614),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_622),
.B(n_610),
.C(n_607),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_644),
.A2(n_641),
.B1(n_616),
.B2(n_623),
.Y(n_664)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_664),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_645),
.B(n_620),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_667),
.B(n_681),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_657),
.A2(n_623),
.B1(n_626),
.B2(n_634),
.Y(n_668)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_668),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_651),
.A2(n_626),
.B1(n_662),
.B2(n_625),
.Y(n_671)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_671),
.Y(n_687)
);

FAx1_ASAP7_75t_SL g672 ( 
.A(n_663),
.B(n_635),
.CI(n_640),
.CON(n_672),
.SN(n_672)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_672),
.B(n_674),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_658),
.B(n_628),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_656),
.A2(n_617),
.B(n_638),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_675),
.A2(n_679),
.B(n_286),
.Y(n_694)
);

XNOR2xp5_ASAP7_75t_L g690 ( 
.A(n_676),
.B(n_678),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_648),
.B(n_632),
.C(n_639),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_SL g695 ( 
.A(n_677),
.B(n_331),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_660),
.A2(n_607),
.B1(n_637),
.B2(n_619),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_SL g681 ( 
.A1(n_643),
.A2(n_585),
.B1(n_469),
.B2(n_316),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_674),
.B(n_654),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_686),
.B(n_691),
.Y(n_702)
);

MAJIxp5_ASAP7_75t_L g688 ( 
.A(n_669),
.B(n_661),
.C(n_649),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_SL g700 ( 
.A(n_688),
.B(n_689),
.Y(n_700)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_669),
.B(n_646),
.C(n_650),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_677),
.B(n_659),
.C(n_642),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_680),
.A2(n_660),
.B(n_340),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_692),
.A2(n_678),
.B(n_672),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_673),
.B(n_354),
.Y(n_693)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_693),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_694),
.B(n_664),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_668),
.B(n_671),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_688),
.Y(n_696)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_696),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_685),
.B(n_666),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_697),
.B(n_704),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_SL g708 ( 
.A1(n_698),
.A2(n_683),
.B(n_684),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_699),
.A2(n_705),
.B(n_682),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_701),
.B(n_690),
.Y(n_709)
);

MAJIxp5_ASAP7_75t_L g704 ( 
.A(n_689),
.B(n_673),
.C(n_665),
.Y(n_704)
);

MAJIxp5_ASAP7_75t_L g705 ( 
.A(n_691),
.B(n_665),
.C(n_670),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_706),
.B(n_709),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_702),
.A2(n_687),
.B(n_692),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_707),
.A2(n_710),
.B(n_672),
.Y(n_715)
);

MAJIxp5_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_698),
.C(n_703),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_700),
.B(n_690),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_714),
.A2(n_715),
.B(n_716),
.Y(n_717)
);

NAND4xp25_ASAP7_75t_L g716 ( 
.A(n_712),
.B(n_670),
.C(n_331),
.D(n_354),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_SL g718 ( 
.A1(n_713),
.A2(n_711),
.B(n_331),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_717),
.B(n_331),
.Y(n_720)
);

MAJIxp5_ASAP7_75t_L g721 ( 
.A(n_720),
.B(n_9),
.C(n_379),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_721),
.B(n_9),
.Y(n_722)
);

XOR2xp5_ASAP7_75t_L g723 ( 
.A(n_722),
.B(n_9),
.Y(n_723)
);


endmodule