module real_jpeg_31988_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_0),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_67),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_0),
.A2(n_67),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_0),
.A2(n_145),
.A3(n_150),
.B1(n_153),
.B2(n_161),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_0),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_0),
.B(n_131),
.Y(n_279)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_1),
.Y(n_339)
);

CKINVDCx11_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_2),
.B(n_503),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B(n_17),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_4),
.Y(n_479)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_6),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_7),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_308)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_7),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_7),
.A2(n_312),
.B1(n_381),
.B2(n_383),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_7),
.A2(n_312),
.B1(n_427),
.B2(n_432),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_7),
.A2(n_312),
.B1(n_470),
.B2(n_475),
.Y(n_469)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_8),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

OAI22x1_ASAP7_75t_SL g28 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_10),
.A2(n_33),
.B1(n_86),
.B2(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_33),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_10),
.A2(n_33),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_12),
.A2(n_342),
.B1(n_343),
.B2(n_345),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_12),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_12),
.A2(n_342),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_12),
.A2(n_342),
.B1(n_457),
.B2(n_460),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_12),
.A2(n_342),
.B1(n_485),
.B2(n_488),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_499),
.B(n_502),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_413),
.B(n_493),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_357),
.B(n_410),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_296),
.Y(n_20)
);

OAI21x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_240),
.B(n_295),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_170),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_23),
.B(n_170),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_104),
.C(n_142),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_24),
.B(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_69),
.B2(n_70),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_71),
.C(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_25),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_25),
.B(n_353),
.C(n_354),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_25),
.B(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_26),
.B(n_401),
.Y(n_400)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_37),
.B1(n_53),
.B2(n_63),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_28),
.A2(n_38),
.B1(n_64),
.B2(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_32),
.Y(n_431)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_36),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_37),
.A2(n_53),
.B(n_63),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_R g481 ( 
.A(n_37),
.B(n_424),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_38),
.B(n_64),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_38),
.A2(n_238),
.B1(n_426),
.B2(n_456),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_53),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_46),
.B2(n_49),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_47),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_52),
.Y(n_160)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_53),
.B(n_67),
.Y(n_265)
);

HB1xp67_ASAP7_75t_SL g424 ( 
.A(n_53),
.Y(n_424)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_56),
.Y(n_166)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_67),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_67),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_67),
.A2(n_197),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_67),
.B(n_247),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_67),
.A2(n_111),
.B(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_68),
.Y(n_462)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_103),
.Y(n_70)
);

OAI211xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_81),
.B(n_84),
.C(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_72),
.B(n_223),
.Y(n_222)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_80),
.B(n_273),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_94),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_82),
.Y(n_203)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_85),
.A2(n_95),
.B1(n_99),
.B2(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_89),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_89),
.Y(n_311)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_93),
.Y(n_258)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_93),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_94),
.A2(n_308),
.B(n_317),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_96),
.B(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_99),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_104),
.A2(n_105),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_104),
.B(n_200),
.C(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_104),
.A2(n_142),
.B1(n_143),
.B2(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_104),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_104),
.B(n_335),
.Y(n_373)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_105),
.Y(n_293)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_122),
.B1(n_131),
.B2(n_132),
.Y(n_105)
);

AOI22x1_ASAP7_75t_L g260 ( 
.A1(n_106),
.A2(n_131),
.B1(n_132),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_106),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_106),
.A2(n_131),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_116),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_107),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_110),
.Y(n_382)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_110),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_111),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_113),
.Y(n_249)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_116),
.B(n_232),
.C(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_116),
.A2(n_235),
.B1(n_380),
.B2(n_387),
.Y(n_379)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_118),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_118),
.Y(n_346)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_123),
.Y(n_261)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_130),
.Y(n_386)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_167),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_144),
.B(n_167),
.Y(n_286)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_168),
.B(n_341),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_169),
.A2(n_308),
.B1(n_336),
.B2(n_340),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_207),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_204),
.B2(n_205),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_172),
.B(n_207),
.C(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_200),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_174),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B(n_188),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_184),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_184),
.Y(n_487)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_200),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_201),
.B(n_279),
.Y(n_280)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_202),
.Y(n_317)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_206),
.B(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_229),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_208),
.B(n_351),
.C(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_208),
.B(n_421),
.C(n_437),
.Y(n_449)
);

MAJx2_ASAP7_75t_L g492 ( 
.A(n_208),
.B(n_449),
.C(n_463),
.Y(n_492)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_209),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_210),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_210),
.A2(n_304),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B(n_218),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_211),
.A2(n_212),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g398 ( 
.A(n_211),
.B(n_323),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_211),
.A2(n_218),
.B(n_469),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_211),
.A2(n_323),
.B1(n_469),
.B2(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_219),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_219),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_221),
.Y(n_488)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_222),
.Y(n_323)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_230),
.B(n_237),
.C(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_231),
.B(n_403),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_236),
.A2(n_237),
.B1(n_259),
.B2(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_236),
.B(n_259),
.C(n_286),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_236),
.A2(n_237),
.B1(n_322),
.B2(n_356),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_237),
.B(n_355),
.C(n_392),
.Y(n_391)
);

AOI21x1_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_289),
.B(n_294),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_283),
.B(n_288),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_266),
.B(n_282),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_262),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_244),
.B(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_259),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_259),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_250),
.B(n_254),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_249),
.Y(n_404)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_259),
.A2(n_270),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_259),
.B(n_307),
.Y(n_351)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_271),
.B(n_281),
.Y(n_266)
);

AOI21x1_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_278),
.B(n_280),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_325),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_300),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_318),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_303),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_329),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_329),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B(n_330),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_352),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_347),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_365),
.C(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_355),
.B(n_422),
.C(n_455),
.Y(n_482)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_356),
.B(n_454),
.Y(n_453)
);

NAND4xp25_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_363),
.D(n_389),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_367),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_372),
.C(n_375),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_375),
.B2(n_376),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_379),
.B2(n_388),
.Y(n_376)
);

OA21x2_ASAP7_75t_SL g440 ( 
.A1(n_377),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_379),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_411),
.B(n_412),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_408),
.B(n_409),
.Y(n_389)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_408),
.C(n_409),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_393),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_399),
.C(n_445),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_398),
.B(n_501),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_406),
.Y(n_399)
);

HB1xp67_ASAP7_75t_SL g418 ( 
.A(n_400),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_401),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_464),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_443),
.B(n_446),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_416),
.B(n_444),
.Y(n_496)
);

XOR2x2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_440),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_438),
.B2(n_439),
.Y(n_417)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_439),
.C(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_423),
.B2(n_437),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B(n_436),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

OAI21x1_ASAP7_75t_SL g495 ( 
.A1(n_446),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_448),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_463),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI221x1_ASAP7_75t_L g493 ( 
.A1(n_464),
.A2(n_466),
.B1(n_494),
.B2(n_495),
.C(n_498),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_489),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_483),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_483),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_480),
.C(n_482),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_480),
.Y(n_491)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx8_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_491),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_500),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_484),
.Y(n_501)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_492),
.Y(n_494)
);


endmodule