module fake_jpeg_29460_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_1),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_62),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_60),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_2),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_2),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_54),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_46),
.B1(n_41),
.B2(n_44),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_69),
.B1(n_4),
.B2(n_5),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_47),
.B1(n_45),
.B2(n_52),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_53),
.B(n_4),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_5),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

OA22x2_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_23),
.B1(n_37),
.B2(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_71),
.B1(n_6),
.B2(n_7),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_11),
.C(n_12),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_103),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.C(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_19),
.B(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_115),
.B(n_118),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_24),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_104),
.C(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_117),
.C(n_116),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_99),
.B1(n_97),
.B2(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_121),
.B1(n_119),
.B2(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_123),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_114),
.B1(n_120),
.B2(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_95),
.C(n_105),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_101),
.A3(n_26),
.B1(n_28),
.B2(n_30),
.C1(n_25),
.C2(n_34),
.Y(n_130)
);


endmodule