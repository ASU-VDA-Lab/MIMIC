module fake_jpeg_19435_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp33_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_54),
.B1(n_50),
.B2(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_94),
.B1(n_86),
.B2(n_62),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_50),
.B1(n_68),
.B2(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_77),
.B1(n_62),
.B2(n_61),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_75),
.B1(n_65),
.B2(n_53),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_92),
.B1(n_90),
.B2(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_96),
.Y(n_108)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_97),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_68),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_69),
.B1(n_74),
.B2(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_80),
.B1(n_67),
.B2(n_78),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_120),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_57),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_56),
.B1(n_66),
.B2(n_60),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_72),
.C(n_71),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_25),
.C(n_43),
.Y(n_139)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_64),
.B1(n_79),
.B2(n_60),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_134),
.B1(n_140),
.B2(n_141),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_142),
.B(n_144),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_29),
.B1(n_49),
.B2(n_47),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_115),
.B1(n_124),
.B2(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_7),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_130),
.B(n_115),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_8),
.B(n_9),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_113),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_11),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_132),
.B1(n_134),
.B2(n_10),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_150),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_153),
.B1(n_147),
.B2(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_159),
.B1(n_152),
.B2(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_154),
.C(n_16),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_14),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_21),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_24),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_32),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_33),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_34),
.B(n_35),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_154),
.C(n_38),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_36),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_40),
.B(n_42),
.Y(n_173)
);


endmodule