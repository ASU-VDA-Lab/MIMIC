module real_aes_831_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g589 ( .A(n_0), .B(n_244), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_1), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g167 ( .A(n_2), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_3), .B(n_526), .Y(n_525) );
NAND2xp33_ASAP7_75t_SL g581 ( .A(n_4), .B(n_184), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_5), .B(n_228), .Y(n_236) );
INVx1_ASAP7_75t_L g574 ( .A(n_6), .Y(n_574) );
INVx1_ASAP7_75t_L g175 ( .A(n_7), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_8), .Y(n_112) );
AOI22xp5_ASAP7_75t_SL g133 ( .A1(n_9), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_9), .Y(n_134) );
OAI22x1_ASAP7_75t_R g136 ( .A1(n_10), .A2(n_80), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_10), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_11), .Y(n_201) );
AND2x2_ASAP7_75t_L g523 ( .A(n_12), .B(n_216), .Y(n_523) );
INVx2_ASAP7_75t_L g157 ( .A(n_13), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g245 ( .A(n_15), .Y(n_245) );
AOI221x1_ASAP7_75t_L g577 ( .A1(n_16), .A2(n_188), .B1(n_528), .B2(n_578), .C(n_580), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_17), .B(n_526), .Y(n_561) );
INVx1_ASAP7_75t_L g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g242 ( .A(n_19), .Y(n_242) );
INVx1_ASAP7_75t_SL g257 ( .A(n_20), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_21), .B(n_178), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_22), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_23), .A2(n_30), .B1(n_514), .B2(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_23), .Y(n_842) );
AOI33xp33_ASAP7_75t_L g282 ( .A1(n_24), .A2(n_54), .A3(n_162), .B1(n_170), .B2(n_283), .B3(n_284), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_25), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_26), .B(n_244), .Y(n_530) );
AOI221xp5_ASAP7_75t_SL g553 ( .A1(n_27), .A2(n_44), .B1(n_526), .B2(n_528), .C(n_554), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_28), .A2(n_829), .B(n_844), .Y(n_828) );
INVx1_ASAP7_75t_L g847 ( .A(n_28), .Y(n_847) );
INVx1_ASAP7_75t_L g193 ( .A(n_29), .Y(n_193) );
NOR3xp33_ASAP7_75t_L g146 ( .A(n_30), .B(n_147), .C(n_338), .Y(n_146) );
INVx1_ASAP7_75t_SL g514 ( .A(n_30), .Y(n_514) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_31), .A2(n_92), .B(n_157), .Y(n_156) );
OR2x2_ASAP7_75t_L g217 ( .A(n_31), .B(n_92), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_32), .B(n_247), .Y(n_565) );
INVxp67_ASAP7_75t_L g576 ( .A(n_33), .Y(n_576) );
AND2x2_ASAP7_75t_L g549 ( .A(n_34), .B(n_215), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_35), .B(n_168), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_36), .A2(n_528), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_37), .B(n_247), .Y(n_555) );
INVx1_ASAP7_75t_L g161 ( .A(n_38), .Y(n_161) );
AND2x2_ASAP7_75t_L g173 ( .A(n_38), .B(n_164), .Y(n_173) );
AND2x2_ASAP7_75t_L g184 ( .A(n_38), .B(n_167), .Y(n_184) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_39), .B(n_111), .C(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g129 ( .A(n_39), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_40), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_41), .B(n_168), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_42), .A2(n_189), .B1(n_224), .B2(n_228), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_43), .B(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_45), .A2(n_84), .B1(n_159), .B2(n_528), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_46), .B(n_178), .Y(n_258) );
INVxp33_ASAP7_75t_L g849 ( .A(n_47), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_48), .B(n_244), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_49), .B(n_155), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_50), .B(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_51), .Y(n_227) );
AND2x2_ASAP7_75t_L g592 ( .A(n_52), .B(n_215), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_53), .B(n_215), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_55), .B(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g166 ( .A(n_56), .Y(n_166) );
INVx1_ASAP7_75t_L g180 ( .A(n_56), .Y(n_180) );
AND2x2_ASAP7_75t_L g214 ( .A(n_57), .B(n_215), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g158 ( .A1(n_58), .A2(n_76), .B1(n_159), .B2(n_168), .C(n_174), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_59), .B(n_168), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_60), .B(n_526), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_61), .B(n_189), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g266 ( .A1(n_62), .A2(n_159), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g540 ( .A(n_63), .B(n_215), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_64), .B(n_247), .Y(n_590) );
INVx1_ASAP7_75t_L g239 ( .A(n_65), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_66), .B(n_244), .Y(n_538) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_67), .B(n_216), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_68), .A2(n_528), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g212 ( .A(n_69), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_70), .B(n_247), .Y(n_531) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_71), .B(n_155), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_72), .A2(n_159), .B(n_211), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_73), .A2(n_133), .B1(n_818), .B2(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g164 ( .A(n_74), .Y(n_164) );
INVx1_ASAP7_75t_L g182 ( .A(n_74), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_75), .B(n_168), .Y(n_285) );
AND2x2_ASAP7_75t_L g259 ( .A(n_77), .B(n_188), .Y(n_259) );
INVx1_ASAP7_75t_L g240 ( .A(n_78), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_79), .A2(n_159), .B(n_256), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_80), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_81), .A2(n_159), .B(n_230), .C(n_234), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_82), .B(n_526), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_83), .A2(n_87), .B1(n_168), .B2(n_526), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_85), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
AND2x2_ASAP7_75t_SL g264 ( .A(n_86), .B(n_188), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_88), .A2(n_159), .B1(n_280), .B2(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_89), .B(n_244), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_90), .B(n_244), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_91), .A2(n_528), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g268 ( .A(n_93), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_94), .B(n_247), .Y(n_537) );
AND2x2_ASAP7_75t_L g286 ( .A(n_95), .B(n_188), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_96), .A2(n_191), .B(n_192), .C(n_195), .Y(n_190) );
INVxp67_ASAP7_75t_L g579 ( .A(n_97), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_98), .B(n_526), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_99), .B(n_247), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_100), .A2(n_528), .B(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_102), .B(n_178), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g839 ( .A1(n_103), .A2(n_840), .B1(n_841), .B2(n_843), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_103), .Y(n_840) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_848), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx8_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx4f_ASAP7_75t_SL g851 ( .A(n_109), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_115), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_114), .B(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_SL g144 ( .A(n_114), .B(n_129), .Y(n_144) );
OR2x6_ASAP7_75t_SL g816 ( .A(n_114), .B(n_128), .Y(n_816) );
OR2x2_ASAP7_75t_L g825 ( .A(n_114), .B(n_129), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_116), .B(n_131), .Y(n_130) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_132), .B1(n_826), .B2(n_828), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
CKINVDCx11_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g827 ( .A(n_120), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp33_ASAP7_75t_L g844 ( .A1(n_124), .A2(n_845), .B(n_846), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g833 ( .A(n_127), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_817), .Y(n_132) );
INVxp33_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B1(n_516), .B2(n_814), .Y(n_140) );
CKINVDCx6p67_ASAP7_75t_R g141 ( .A(n_142), .Y(n_141) );
CKINVDCx11_ASAP7_75t_R g821 ( .A(n_142), .Y(n_821) );
INVx3_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_144), .Y(n_143) );
AOI211xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_409), .B(n_512), .C(n_515), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_146), .A2(n_409), .B(n_512), .Y(n_819) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_148), .A2(n_410), .B(n_514), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_148), .B(n_487), .Y(n_837) );
NOR2x1_ASAP7_75t_L g148 ( .A(n_149), .B(n_316), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_299), .Y(n_149) );
AOI221xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_218), .B1(n_260), .B2(n_274), .C(n_289), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_205), .Y(n_151) );
NAND2x1_ASAP7_75t_SL g325 ( .A(n_152), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g352 ( .A(n_152), .B(n_322), .Y(n_352) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_152), .Y(n_398) );
AND2x2_ASAP7_75t_L g406 ( .A(n_152), .B(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g510 ( .A(n_152), .Y(n_510) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_186), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_154), .Y(n_288) );
INVx1_ASAP7_75t_L g304 ( .A(n_154), .Y(n_304) );
AND2x4_ASAP7_75t_L g311 ( .A(n_154), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g321 ( .A(n_154), .B(n_186), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_154), .B(n_307), .Y(n_348) );
INVx1_ASAP7_75t_L g359 ( .A(n_154), .Y(n_359) );
INVxp67_ASAP7_75t_L g393 ( .A(n_154), .Y(n_393) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_185), .Y(n_154) );
INVx2_ASAP7_75t_SL g234 ( .A(n_155), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_155), .A2(n_561), .B(n_562), .Y(n_560) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_157), .B(n_217), .Y(n_216) );
AND2x4_ASAP7_75t_L g228 ( .A(n_157), .B(n_217), .Y(n_228) );
INVxp67_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_159), .A2(n_168), .B1(n_573), .B2(n_575), .Y(n_572) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_165), .Y(n_159) );
NOR2x1p5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx1_ASAP7_75t_L g284 ( .A(n_162), .Y(n_284) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x6_ASAP7_75t_L g176 ( .A(n_163), .B(n_170), .Y(n_176) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x6_ASAP7_75t_L g244 ( .A(n_164), .B(n_179), .Y(n_244) );
AND2x6_ASAP7_75t_L g528 ( .A(n_165), .B(n_173), .Y(n_528) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g170 ( .A(n_166), .Y(n_170) );
AND2x4_ASAP7_75t_L g247 ( .A(n_166), .B(n_181), .Y(n_247) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
INVx1_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_172), .Y(n_168) );
INVx1_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVxp33_ASAP7_75t_L g283 ( .A(n_170), .Y(n_283) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
INVxp67_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_176), .A2(n_183), .B(n_212), .C(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g233 ( .A(n_176), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_176), .A2(n_194), .B1(n_239), .B2(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_176), .A2(n_183), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_176), .A2(n_183), .B(n_268), .C(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
AND2x4_ASAP7_75t_L g526 ( .A(n_178), .B(n_184), .Y(n_526) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_183), .A2(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_183), .B(n_228), .Y(n_248) );
INVx1_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_183), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_183), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_183), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_183), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_183), .A2(n_564), .B(n_565), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_183), .A2(n_589), .B(n_590), .Y(n_588) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_184), .Y(n_195) );
INVx2_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_186), .B(n_207), .Y(n_292) );
INVx1_ASAP7_75t_L g310 ( .A(n_186), .Y(n_310) );
INVx1_ASAP7_75t_L g357 ( .A(n_186), .Y(n_357) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_198), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B1(n_196), .B2(n_197), .Y(n_187) );
INVx3_ASAP7_75t_L g197 ( .A(n_188), .Y(n_197) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_189), .B(n_200), .Y(n_199) );
AOI21x1_ASAP7_75t_L g585 ( .A1(n_189), .A2(n_586), .B(n_592), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_194), .B(n_228), .C(n_581), .Y(n_580) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_197), .A2(n_208), .B(n_214), .Y(n_207) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_197), .A2(n_208), .B(n_214), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_205), .B(n_329), .Y(n_334) );
AND2x2_ASAP7_75t_L g346 ( .A(n_205), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g365 ( .A(n_205), .B(n_311), .Y(n_365) );
INVx1_ASAP7_75t_L g374 ( .A(n_205), .Y(n_374) );
AND2x2_ASAP7_75t_L g422 ( .A(n_205), .B(n_321), .Y(n_422) );
OR2x2_ASAP7_75t_L g465 ( .A(n_205), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_L g305 ( .A(n_206), .B(n_306), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_206), .B(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g287 ( .A(n_207), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_207), .B(n_307), .Y(n_385) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_207), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_215), .Y(n_252) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_215), .A2(n_553), .B(n_557), .Y(n_552) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_249), .Y(n_219) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_220), .B(n_344), .Y(n_389) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g351 ( .A(n_221), .B(n_342), .Y(n_351) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
INVx1_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
AND2x4_ASAP7_75t_L g297 ( .A(n_222), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g301 ( .A(n_222), .Y(n_301) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_222), .Y(n_337) );
AND2x2_ASAP7_75t_L g507 ( .A(n_222), .B(n_263), .Y(n_507) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .C(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_228), .A2(n_266), .B(n_270), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_228), .A2(n_525), .B(n_527), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_228), .B(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_228), .B(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_228), .B(n_579), .Y(n_578) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_234), .A2(n_278), .B(n_286), .Y(n_277) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_234), .A2(n_278), .B(n_286), .Y(n_307) );
AOI21x1_ASAP7_75t_L g600 ( .A1(n_234), .A2(n_601), .B(n_604), .Y(n_600) );
INVx3_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
INVx2_ASAP7_75t_L g315 ( .A(n_235), .Y(n_315) );
NOR2x1_ASAP7_75t_SL g332 ( .A(n_235), .B(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g370 ( .A(n_235), .B(n_251), .Y(n_370) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_241), .B(n_248), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B1(n_245), .B2(n_246), .Y(n_241) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g444 ( .A(n_249), .Y(n_444) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
INVx1_ASAP7_75t_L g342 ( .A(n_251), .Y(n_342) );
INVx1_ASAP7_75t_L g402 ( .A(n_251), .Y(n_402) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_251), .Y(n_421) );
OR2x2_ASAP7_75t_L g427 ( .A(n_251), .B(n_263), .Y(n_427) );
AND2x2_ASAP7_75t_L g471 ( .A(n_251), .B(n_298), .Y(n_471) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_259), .Y(n_251) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_252), .A2(n_534), .B(n_540), .Y(n_533) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_252), .A2(n_543), .B(n_549), .Y(n_542) );
AO21x2_ASAP7_75t_L g681 ( .A1(n_252), .A2(n_543), .B(n_549), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_272), .Y(n_261) );
AND2x2_ASAP7_75t_L g313 ( .A(n_262), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g467 ( .A(n_262), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g472 ( .A(n_262), .Y(n_472) );
AND2x2_ASAP7_75t_L g484 ( .A(n_262), .B(n_370), .Y(n_484) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_271), .Y(n_262) );
INVx4_ASAP7_75t_L g295 ( .A(n_263), .Y(n_295) );
INVx2_ASAP7_75t_L g345 ( .A(n_263), .Y(n_345) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_263), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_263), .B(n_403), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_263), .B(n_273), .Y(n_476) );
AND2x2_ASAP7_75t_L g502 ( .A(n_263), .B(n_315), .Y(n_502) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x4_ASAP7_75t_L g404 ( .A(n_271), .B(n_295), .Y(n_404) );
AND2x2_ASAP7_75t_L g331 ( .A(n_272), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g349 ( .A(n_272), .B(n_336), .Y(n_349) );
INVx1_ASAP7_75t_L g383 ( .A(n_272), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_272), .B(n_297), .Y(n_439) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_273), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_274), .A2(n_356), .B1(n_500), .B2(n_503), .Y(n_499) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_287), .Y(n_274) );
INVx1_ASAP7_75t_L g429 ( .A(n_275), .Y(n_429) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g452 ( .A(n_276), .B(n_324), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_276), .B(n_324), .Y(n_461) );
INVx2_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x4_ASAP7_75t_L g322 ( .A(n_277), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_277), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_279), .B(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_288), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_291), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g396 ( .A(n_291), .B(n_311), .Y(n_396) );
INVx2_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g434 ( .A(n_292), .B(n_348), .Y(n_434) );
INVxp33_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g415 ( .A(n_294), .Y(n_415) );
NOR2x1_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x4_ASAP7_75t_SL g336 ( .A(n_295), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
INVx2_ASAP7_75t_L g425 ( .A(n_296), .Y(n_425) );
NAND2xp33_ASAP7_75t_SL g500 ( .A(n_296), .B(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g366 ( .A(n_297), .B(n_345), .Y(n_366) );
AND2x2_ASAP7_75t_L g300 ( .A(n_298), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g403 ( .A(n_298), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_302), .B1(n_308), .B2(n_313), .Y(n_299) );
AND2x2_ASAP7_75t_L g328 ( .A(n_300), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g433 ( .A(n_300), .Y(n_433) );
INVx1_ASAP7_75t_L g382 ( .A(n_301), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_302), .A2(n_341), .B1(n_346), .B2(n_349), .Y(n_340) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_L g466 ( .A(n_303), .Y(n_466) );
BUFx3_ASAP7_75t_L g431 ( .A(n_304), .Y(n_431) );
INVx1_ASAP7_75t_L g454 ( .A(n_305), .Y(n_454) );
AND2x2_ASAP7_75t_L g392 ( .A(n_306), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g459 ( .A(n_306), .B(n_324), .Y(n_459) );
INVx1_ASAP7_75t_L g493 ( .A(n_306), .Y(n_493) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI21xp33_ASAP7_75t_L g330 ( .A1(n_308), .A2(n_331), .B(n_333), .Y(n_330) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_308), .A2(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g441 ( .A(n_310), .Y(n_441) );
AND2x2_ASAP7_75t_L g458 ( .A(n_310), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g448 ( .A(n_311), .B(n_407), .Y(n_448) );
AND2x2_ASAP7_75t_L g451 ( .A(n_311), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g460 ( .A(n_311), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g405 ( .A(n_314), .B(n_404), .Y(n_405) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_315), .B(n_344), .Y(n_343) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_315), .B(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_327), .B(n_330), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_325), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_320), .A2(n_336), .B1(n_361), .B2(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_324), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_326), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_326), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g468 ( .A(n_329), .Y(n_468) );
AND2x2_ASAP7_75t_L g455 ( .A(n_332), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_R g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_336), .B(n_419), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_338), .Y(n_513) );
OR3x2_ASAP7_75t_L g836 ( .A(n_338), .B(n_411), .C(n_837), .Y(n_836) );
NAND3x1_ASAP7_75t_SL g338 ( .A(n_339), .B(n_353), .C(n_367), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_350), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_341), .A2(n_451), .B1(n_453), .B2(n_455), .Y(n_450) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_342), .B(n_381), .Y(n_395) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_347), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g416 ( .A(n_347), .B(n_357), .Y(n_416) );
AND2x2_ASAP7_75t_L g440 ( .A(n_347), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_351), .A2(n_447), .B(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_L g498 ( .A(n_351), .B(n_377), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_352), .A2(n_505), .B1(n_508), .B2(n_511), .Y(n_504) );
AOI21xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_360), .B(n_364), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
BUFx2_ASAP7_75t_L g474 ( .A(n_357), .Y(n_474) );
INVx1_ASAP7_75t_SL g481 ( .A(n_357), .Y(n_481) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_358), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_387), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g376 ( .A(n_370), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_370), .B(n_381), .Y(n_462) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_378), .B(n_384), .Y(n_375) );
OR2x6_ASAP7_75t_L g432 ( .A(n_377), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
OR2x2_ASAP7_75t_L g509 ( .A(n_385), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_386), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_397), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_394), .B2(n_396), .Y(n_388) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_391), .Y(n_489) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_405), .B2(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_485), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_435), .C(n_463), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_423), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_417), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g456 ( .A(n_420), .Y(n_456) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_428), .B1(n_432), .B2(n_434), .Y(n_423) );
NAND2x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_425), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_427), .B(n_433), .Y(n_503) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx3_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
INVx2_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_449), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_437), .B(n_446), .Y(n_436) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_440), .B1(n_442), .B2(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_445), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_450), .B(n_457), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_452), .B(n_493), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B(n_462), .Y(n_457) );
INVx1_ASAP7_75t_L g477 ( .A(n_460), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B(n_469), .C(n_478), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_466), .A2(n_497), .B(n_499), .C(n_504), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B1(n_475), .B2(n_477), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVxp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_SL g512 ( .A1(n_485), .A2(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
AOI21xp33_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_490), .B(n_494), .Y(n_488) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVxp33_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_515), .B(n_821), .Y(n_820) );
AO22x2_ASAP7_75t_L g818 ( .A1(n_516), .A2(n_815), .B1(n_819), .B2(n_820), .Y(n_818) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_725), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_647), .C(n_697), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_614), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_550), .B1(n_567), .B2(n_597), .C(n_606), .Y(n_520) );
INVx1_ASAP7_75t_SL g696 ( .A(n_521), .Y(n_696) );
AND2x4_ASAP7_75t_SL g521 ( .A(n_522), .B(n_532), .Y(n_521) );
INVx2_ASAP7_75t_L g618 ( .A(n_522), .Y(n_618) );
OR2x2_ASAP7_75t_L g640 ( .A(n_522), .B(n_631), .Y(n_640) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_522), .Y(n_655) );
INVx5_ASAP7_75t_L g662 ( .A(n_522), .Y(n_662) );
AND2x4_ASAP7_75t_L g668 ( .A(n_522), .B(n_542), .Y(n_668) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_522), .B(n_599), .Y(n_671) );
OR2x2_ASAP7_75t_L g680 ( .A(n_522), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g687 ( .A(n_522), .B(n_533), .Y(n_687) );
AND2x2_ASAP7_75t_L g788 ( .A(n_522), .B(n_541), .Y(n_788) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx3_ASAP7_75t_SL g639 ( .A(n_532), .Y(n_639) );
AND2x2_ASAP7_75t_L g683 ( .A(n_532), .B(n_599), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_532), .A2(n_687), .B(n_688), .Y(n_686) );
AND2x2_ASAP7_75t_L g724 ( .A(n_532), .B(n_662), .Y(n_724) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_541), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_533), .B(n_542), .Y(n_605) );
OR2x2_ASAP7_75t_L g609 ( .A(n_533), .B(n_542), .Y(n_609) );
INVx1_ASAP7_75t_L g617 ( .A(n_533), .Y(n_617) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_533), .Y(n_629) );
INVx2_ASAP7_75t_L g637 ( .A(n_533), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_533), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g746 ( .A(n_533), .B(n_631), .Y(n_746) );
AND2x2_ASAP7_75t_L g761 ( .A(n_533), .B(n_599), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g630 ( .A(n_542), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_542), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_550), .B(n_754), .Y(n_753) );
NOR2x1p5_ASAP7_75t_L g550 ( .A(n_551), .B(n_558), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g583 ( .A(n_552), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_552), .B(n_559), .Y(n_612) );
INVx1_ASAP7_75t_L g622 ( .A(n_552), .Y(n_622) );
INVx2_ASAP7_75t_L g645 ( .A(n_552), .Y(n_645) );
INVx2_ASAP7_75t_L g651 ( .A(n_552), .Y(n_651) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_552), .Y(n_721) );
OR2x2_ASAP7_75t_L g752 ( .A(n_552), .B(n_559), .Y(n_752) );
OR2x2_ASAP7_75t_L g768 ( .A(n_558), .B(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_SL g570 ( .A(n_559), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g595 ( .A(n_559), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g632 ( .A(n_559), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g644 ( .A(n_559), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g657 ( .A(n_559), .B(n_623), .Y(n_657) );
OR2x2_ASAP7_75t_L g665 ( .A(n_559), .B(n_571), .Y(n_665) );
INVx2_ASAP7_75t_L g692 ( .A(n_559), .Y(n_692) );
INVx1_ASAP7_75t_L g710 ( .A(n_559), .Y(n_710) );
NOR2xp33_ASAP7_75t_R g743 ( .A(n_559), .B(n_584), .Y(n_743) );
OR2x6_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_568), .B(n_593), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_568), .A2(n_635), .B1(n_638), .B2(n_641), .Y(n_634) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_582), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g649 ( .A(n_570), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g684 ( .A(n_570), .B(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_L g763 ( .A(n_570), .B(n_741), .Y(n_763) );
INVx3_ASAP7_75t_L g596 ( .A(n_571), .Y(n_596) );
AND2x4_ASAP7_75t_L g623 ( .A(n_571), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_571), .B(n_584), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_571), .B(n_645), .Y(n_690) );
AND2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_692), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_571), .B(n_583), .Y(n_732) );
INVx1_ASAP7_75t_L g802 ( .A(n_571), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_571), .B(n_720), .Y(n_813) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g594 ( .A(n_584), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_584), .B(n_596), .Y(n_613) );
INVx2_ASAP7_75t_L g624 ( .A(n_584), .Y(n_624) );
AND2x2_ASAP7_75t_L g650 ( .A(n_584), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g666 ( .A(n_584), .B(n_645), .Y(n_666) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_584), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_584), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g755 ( .A(n_584), .Y(n_755) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_591), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_594), .B(n_622), .Y(n_633) );
AOI221x1_ASAP7_75t_SL g727 ( .A1(n_595), .A2(n_728), .B1(n_731), .B2(n_733), .C(n_737), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_595), .B(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g785 ( .A(n_595), .B(n_650), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_595), .B(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g716 ( .A(n_596), .B(n_644), .Y(n_716) );
AND2x2_ASAP7_75t_L g754 ( .A(n_596), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_605), .Y(n_598) );
AND2x2_ASAP7_75t_L g607 ( .A(n_599), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g702 ( .A(n_599), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_599), .B(n_618), .Y(n_707) );
AND2x4_ASAP7_75t_L g736 ( .A(n_599), .B(n_637), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_599), .B(n_668), .Y(n_772) );
OR2x2_ASAP7_75t_L g790 ( .A(n_599), .B(n_721), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_599), .B(n_681), .Y(n_800) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g631 ( .A(n_600), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g656 ( .A(n_605), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_605), .A2(n_664), .B1(n_667), .B2(n_669), .Y(n_663) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
INVx2_ASAP7_75t_L g619 ( .A(n_607), .Y(n_619) );
AND2x2_ASAP7_75t_L g758 ( .A(n_608), .B(n_618), .Y(n_758) );
AND2x2_ASAP7_75t_L g804 ( .A(n_608), .B(n_671), .Y(n_804) );
AND2x2_ASAP7_75t_L g809 ( .A(n_608), .B(n_660), .Y(n_809) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g778 ( .A1(n_610), .A2(n_680), .A3(n_760), .B1(n_779), .B2(n_781), .Y(n_778) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g646 ( .A(n_613), .Y(n_646) );
AOI211xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_620), .B(n_625), .C(n_634), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_617), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_618), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g798 ( .A(n_618), .Y(n_798) );
AND2x2_ASAP7_75t_L g708 ( .A(n_620), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_621), .B(n_623), .Y(n_620) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_621), .Y(n_808) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_622), .Y(n_677) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_622), .Y(n_777) );
INVx1_ASAP7_75t_L g674 ( .A(n_623), .Y(n_674) );
AND2x2_ASAP7_75t_L g740 ( .A(n_623), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_623), .B(n_751), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_632), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_627), .A2(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_SL g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g636 ( .A(n_631), .B(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g660 ( .A(n_631), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_636), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g767 ( .A(n_636), .Y(n_767) );
AND2x2_ASAP7_75t_L g797 ( .A(n_636), .B(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_637), .Y(n_774) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_639), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g714 ( .A(n_640), .Y(n_714) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g673 ( .A(n_644), .B(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_645), .Y(n_741) );
AND2x2_ASAP7_75t_L g750 ( .A(n_646), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_670), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B1(n_657), .B2(n_658), .C(n_663), .Y(n_648) );
INVx1_ASAP7_75t_L g769 ( .A(n_650), .Y(n_769) );
INVxp33_ASAP7_75t_SL g801 ( .A(n_650), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_652), .A2(n_748), .B(n_756), .Y(n_747) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_656), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g669 ( .A(n_657), .Y(n_669) );
AND2x2_ASAP7_75t_L g704 ( .A(n_657), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g723 ( .A(n_657), .B(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_657), .A2(n_785), .B1(n_786), .B2(n_789), .Y(n_784) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
OR2x2_ASAP7_75t_L g679 ( .A(n_660), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_660), .B(n_668), .Y(n_718) );
AND2x4_ASAP7_75t_L g735 ( .A(n_662), .B(n_681), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_662), .B(n_736), .Y(n_782) );
AND2x2_ASAP7_75t_L g794 ( .A(n_662), .B(n_746), .Y(n_794) );
NAND2xp33_ASAP7_75t_L g779 ( .A(n_664), .B(n_780), .Y(n_779) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_SL g722 ( .A(n_665), .Y(n_722) );
INVx1_ASAP7_75t_L g793 ( .A(n_666), .Y(n_793) );
INVx2_ASAP7_75t_SL g745 ( .A(n_668), .Y(n_745) );
AOI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_672), .B(n_675), .C(n_693), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B(n_682), .C(n_686), .Y(n_675) );
OR2x6_ASAP7_75t_SL g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g705 ( .A(n_677), .Y(n_705) );
INVx1_ASAP7_75t_SL g730 ( .A(n_680), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_680), .B(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_685), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g771 ( .A1(n_689), .A2(n_772), .B1(n_773), .B2(n_775), .Y(n_771) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_703), .B(n_706), .C(n_711), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_723), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g803 ( .A1(n_722), .A2(n_804), .B1(n_805), .B2(n_809), .C1(n_810), .C2(n_812), .Y(n_803) );
INVx2_ASAP7_75t_L g738 ( .A(n_724), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_764), .C(n_783), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_747), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_735), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_736), .B(n_798), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_742), .B2(n_744), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVxp33_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_745), .B(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_753), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_753), .A2(n_757), .B1(n_759), .B2(n_762), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
CKINVDCx16_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
OAI211xp5_ASAP7_75t_SL g764 ( .A1(n_765), .A2(n_768), .B(n_770), .C(n_778), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_791), .C(n_803), .Y(n_783) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_795), .B(n_802), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_799), .B(n_801), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
INVx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_831), .B(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_833), .Y(n_832) );
INVxp67_ASAP7_75t_L g845 ( .A(n_834), .Y(n_845) );
AOI22x1_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B1(n_838), .B2(n_839), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g843 ( .A(n_841), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
endmodule