module fake_netlist_1_5541_n_473 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_473);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_473;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g67 ( .A(n_34), .B(n_21), .Y(n_67) );
BUFx6f_ASAP7_75t_L g68 ( .A(n_11), .Y(n_68) );
INVxp67_ASAP7_75t_SL g69 ( .A(n_22), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_53), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_20), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_5), .Y(n_72) );
INVxp33_ASAP7_75t_SL g73 ( .A(n_32), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_58), .Y(n_74) );
BUFx3_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_25), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_55), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_50), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_59), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_52), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_40), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_62), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_9), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_44), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_57), .Y(n_88) );
BUFx8_ASAP7_75t_SL g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_19), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_26), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_0), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_16), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_39), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_10), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_61), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_42), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_27), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_102), .B(n_0), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_75), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_75), .B(n_1), .Y(n_106) );
CKINVDCx6p67_ASAP7_75t_R g107 ( .A(n_98), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
INVx3_ASAP7_75t_L g109 ( .A(n_68), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_102), .B(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
OR2x6_ASAP7_75t_L g118 ( .A(n_72), .B(n_31), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_72), .B(n_2), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_91), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_68), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_91), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_68), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_78), .A2(n_33), .B(n_66), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_68), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_105), .B(n_98), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
NAND3x1_ASAP7_75t_L g130 ( .A(n_119), .B(n_99), .C(n_94), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_107), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
BUFx4f_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_107), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
INVx5_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_107), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_105), .A2(n_93), .B1(n_88), .B2(n_83), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_125), .B(n_79), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_105), .B(n_93), .Y(n_143) );
OR2x6_ASAP7_75t_L g144 ( .A(n_118), .B(n_85), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_108), .B(n_84), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_118), .A2(n_117), .B1(n_112), .B2(n_115), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
INVx2_ASAP7_75t_SL g149 ( .A(n_136), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_128), .B(n_108), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_143), .B(n_112), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_136), .A2(n_118), .B1(n_119), .B2(n_117), .Y(n_156) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
OR2x4_ASAP7_75t_L g161 ( .A(n_133), .B(n_104), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_144), .A2(n_121), .B1(n_115), .B2(n_116), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_144), .B(n_104), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_130), .A2(n_121), .B1(n_116), .B2(n_73), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_145), .B(n_70), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_139), .B(n_95), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_141), .B(n_96), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_144), .A2(n_94), .B1(n_85), .B2(n_90), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_139), .B(n_103), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_139), .B(n_69), .Y(n_181) );
BUFx12f_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_151), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_167), .B(n_139), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_157), .A2(n_136), .B1(n_146), .B2(n_139), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_173), .A2(n_139), .B1(n_141), .B2(n_142), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
AOI33xp33_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_90), .A3(n_99), .B1(n_92), .B2(n_80), .B3(n_81), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_167), .B(n_92), .Y(n_190) );
INVxp67_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_157), .A2(n_130), .B1(n_142), .B2(n_76), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_157), .B(n_68), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_152), .B(n_100), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_173), .A2(n_68), .B1(n_97), .B2(n_86), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_167), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_150), .B(n_89), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_167), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_172), .B(n_79), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_176), .B(n_3), .Y(n_208) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_156), .A2(n_81), .B(n_80), .Y(n_209) );
HAxp5_ASAP7_75t_L g210 ( .A(n_176), .B(n_161), .CON(n_210), .SN(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_149), .B(n_82), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_164), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_206), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_187), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_193), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_173), .B1(n_177), .B2(n_162), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_189), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_191), .B(n_161), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_201), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_182), .A2(n_149), .B1(n_170), .B2(n_164), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_188), .B(n_161), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_210), .B(n_153), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g228 ( .A1(n_183), .A2(n_163), .B1(n_153), .B2(n_168), .Y(n_228) );
OAI21xp33_ASAP7_75t_SL g229 ( .A1(n_198), .A2(n_165), .B(n_170), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_208), .B(n_165), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_197), .A2(n_168), .B1(n_169), .B2(n_158), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_207), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_197), .A2(n_168), .B1(n_169), .B2(n_158), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_207), .A2(n_180), .B(n_169), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_197), .A2(n_154), .B1(n_171), .B2(n_178), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_214), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_214), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_208), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_200), .B(n_202), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_200), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_240), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_227), .A2(n_190), .B1(n_197), .B2(n_199), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_227), .A2(n_239), .B1(n_190), .B2(n_228), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
AOI221xp5_ASAP7_75t_SL g247 ( .A1(n_229), .A2(n_205), .B1(n_196), .B2(n_195), .C(n_194), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_226), .A2(n_190), .B1(n_192), .B2(n_213), .C(n_202), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_241), .A2(n_201), .B1(n_203), .B2(n_190), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_231), .A2(n_213), .B1(n_192), .B2(n_203), .Y(n_253) );
AOI222xp33_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_210), .B1(n_185), .B2(n_201), .C1(n_154), .C2(n_189), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_213), .B1(n_201), .B2(n_189), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_229), .A2(n_213), .B1(n_174), .B2(n_206), .C(n_210), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_238), .A2(n_201), .B1(n_189), .B2(n_209), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_234), .A2(n_212), .B(n_211), .Y(n_259) );
NAND3xp33_ASAP7_75t_L g260 ( .A(n_234), .B(n_204), .C(n_126), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_218), .B(n_189), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_222), .A2(n_209), .B1(n_184), .B2(n_212), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g264 ( .A(n_247), .B(n_232), .C(n_237), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_243), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_209), .B1(n_221), .B2(n_237), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_242), .A2(n_238), .B1(n_222), .B2(n_223), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_251), .B(n_223), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_254), .A2(n_233), .B1(n_219), .B2(n_225), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_252), .B(n_233), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_253), .A2(n_236), .B1(n_184), .B2(n_224), .Y(n_272) );
OAI31xp33_ASAP7_75t_L g273 ( .A1(n_242), .A2(n_236), .A3(n_184), .B(n_230), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_235), .B(n_179), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_252), .B(n_220), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_254), .A2(n_184), .B1(n_220), .B2(n_211), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_243), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_249), .A2(n_220), .B1(n_212), .B2(n_211), .Y(n_279) );
OAI33xp33_ASAP7_75t_L g280 ( .A1(n_251), .A2(n_82), .A3(n_101), .B1(n_87), .B2(n_86), .B3(n_77), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_256), .A2(n_87), .B1(n_101), .B2(n_77), .C(n_181), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_246), .B(n_125), .Y(n_282) );
OAI33xp33_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_113), .A3(n_178), .B1(n_179), .B2(n_7), .B3(n_8), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_258), .B(n_261), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_246), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_268), .B(n_246), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_268), .B(n_248), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_265), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
AOI33xp33_ASAP7_75t_L g290 ( .A1(n_266), .A2(n_244), .A3(n_263), .B1(n_261), .B2(n_257), .B3(n_250), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_277), .B(n_248), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_278), .B(n_259), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
AND2x4_ASAP7_75t_SL g294 ( .A(n_271), .B(n_248), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_274), .A2(n_260), .B(n_259), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_265), .Y(n_297) );
OAI31xp33_ASAP7_75t_L g298 ( .A1(n_273), .A2(n_260), .A3(n_255), .B(n_262), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_285), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_278), .B(n_262), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_277), .B(n_125), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_264), .A2(n_67), .B(n_211), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
AOI31xp33_ASAP7_75t_L g304 ( .A1(n_276), .A2(n_4), .A3(n_5), .B(n_6), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_265), .A2(n_125), .B(n_204), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_270), .A2(n_212), .B1(n_204), .B2(n_125), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_271), .B(n_113), .Y(n_308) );
OAI33xp33_ASAP7_75t_L g309 ( .A1(n_267), .A2(n_113), .A3(n_6), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_309) );
NOR2xp33_ASAP7_75t_SL g310 ( .A(n_273), .B(n_204), .Y(n_310) );
NAND4xp25_ASAP7_75t_L g311 ( .A(n_281), .B(n_109), .C(n_122), .D(n_113), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_264), .B(n_51), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_275), .B(n_124), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_269), .B(n_4), .Y(n_315) );
AND3x2_ASAP7_75t_L g316 ( .A(n_310), .B(n_281), .C(n_275), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_306), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_314), .B(n_269), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_289), .B(n_274), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_288), .B(n_282), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_314), .B(n_279), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_289), .B(n_272), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_308), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_308), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_308), .Y(n_327) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_294), .B(n_282), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_289), .B(n_272), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_294), .B(n_12), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_288), .B(n_126), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_124), .Y(n_332) );
OAI31xp33_ASAP7_75t_L g333 ( .A1(n_315), .A2(n_122), .A3(n_109), .B(n_283), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_304), .A2(n_280), .B1(n_204), .B2(n_15), .Y(n_334) );
OAI33xp33_ASAP7_75t_L g335 ( .A1(n_311), .A2(n_13), .A3(n_14), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_124), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_286), .B(n_14), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_287), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_287), .B(n_124), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_291), .B(n_124), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_291), .B(n_124), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_310), .A2(n_280), .B(n_175), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_290), .B(n_17), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_309), .B(n_313), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_309), .A2(n_122), .B1(n_124), .B2(n_126), .C(n_110), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_322), .B(n_324), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_338), .B(n_299), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_328), .B(n_288), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_328), .B(n_297), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_339), .B(n_303), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_334), .A2(n_298), .B(n_312), .Y(n_360) );
AND4x1_ASAP7_75t_L g361 ( .A(n_335), .B(n_302), .C(n_307), .D(n_305), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_343), .B(n_297), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_318), .B(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_325), .B(n_297), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_344), .A2(n_292), .B1(n_296), .B2(n_293), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_349), .B(n_307), .C(n_126), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_326), .B(n_292), .Y(n_369) );
XNOR2xp5_ASAP7_75t_L g370 ( .A(n_316), .B(n_292), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_345), .B(n_293), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_327), .B(n_293), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_321), .B(n_293), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_330), .B(n_296), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_341), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_350), .B(n_126), .C(n_111), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_350), .A2(n_126), .B1(n_111), .B2(n_114), .C(n_120), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g380 ( .A1(n_337), .A2(n_296), .B(n_301), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_347), .B(n_296), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_351), .B(n_123), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_305), .B1(n_123), .B2(n_120), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_353), .A2(n_110), .B(n_111), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_329), .B(n_123), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_342), .B(n_123), .Y(n_386) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_348), .B(n_120), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_345), .A2(n_110), .B(n_111), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_331), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_323), .B(n_120), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_364), .B(n_319), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_370), .A2(n_333), .B(n_320), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_360), .A2(n_346), .B(n_331), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_391), .Y(n_401) );
AOI211x1_ASAP7_75t_L g402 ( .A1(n_361), .A2(n_336), .B(n_114), .C(n_111), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_375), .B(n_114), .Y(n_403) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_357), .B(n_148), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_387), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_387), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_385), .B(n_23), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_376), .B(n_29), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_380), .B(n_148), .Y(n_410) );
AOI32xp33_ASAP7_75t_L g411 ( .A1(n_367), .A2(n_30), .A3(n_35), .B1(n_36), .B2(n_37), .Y(n_411) );
XOR2x1_ASAP7_75t_L g412 ( .A(n_365), .B(n_38), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_376), .B(n_41), .Y(n_413) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_390), .Y(n_414) );
XNOR2x2_ASAP7_75t_L g415 ( .A(n_378), .B(n_43), .Y(n_415) );
INVxp33_ASAP7_75t_L g416 ( .A(n_372), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_390), .Y(n_418) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_368), .B(n_45), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_381), .B(n_46), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_355), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_373), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_366), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
XOR2xp5_ASAP7_75t_L g425 ( .A(n_377), .B(n_47), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_148), .B(n_134), .C(n_127), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_384), .A2(n_48), .B(n_49), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_371), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_362), .B(n_54), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
INVxp33_ASAP7_75t_SL g431 ( .A(n_386), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_389), .B(n_56), .Y(n_432) );
XNOR2xp5_ASAP7_75t_L g433 ( .A(n_371), .B(n_63), .Y(n_433) );
XNOR2x2_ASAP7_75t_L g434 ( .A(n_383), .B(n_64), .Y(n_434) );
AO22x2_ASAP7_75t_L g435 ( .A1(n_388), .A2(n_127), .B1(n_134), .B2(n_391), .Y(n_435) );
XOR2xp5_ASAP7_75t_L g436 ( .A(n_370), .B(n_127), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_356), .Y(n_437) );
XOR2x2_ASAP7_75t_L g438 ( .A(n_370), .B(n_127), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_370), .B(n_134), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_363), .B(n_134), .Y(n_440) );
AO21x1_ASAP7_75t_L g441 ( .A1(n_387), .A2(n_360), .B(n_380), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_391), .B(n_390), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_414), .B(n_418), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_423), .A2(n_397), .B1(n_437), .B2(n_406), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_403), .A2(n_436), .B(n_441), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_442), .B(n_437), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_405), .A2(n_399), .B(n_400), .Y(n_448) );
AOI322xp5_ASAP7_75t_L g449 ( .A1(n_396), .A2(n_421), .A3(n_398), .B1(n_408), .B2(n_393), .C1(n_424), .C2(n_422), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_404), .A2(n_410), .B(n_399), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_439), .A2(n_431), .B1(n_433), .B2(n_416), .Y(n_451) );
OAI211xp5_ASAP7_75t_SL g452 ( .A1(n_411), .A2(n_394), .B(n_428), .C(n_413), .Y(n_452) );
OAI222xp33_ASAP7_75t_R g453 ( .A1(n_434), .A2(n_425), .B1(n_417), .B2(n_430), .C1(n_415), .C2(n_401), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_448), .A2(n_438), .B1(n_409), .B2(n_429), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_445), .A2(n_426), .B(n_440), .C(n_420), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_444), .A2(n_435), .B1(n_402), .B2(n_419), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_452), .B(n_420), .C(n_432), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_450), .B(n_427), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_449), .A2(n_412), .B(n_427), .C(n_407), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_460), .A2(n_451), .B(n_443), .Y(n_461) );
XNOR2xp5_ASAP7_75t_L g462 ( .A(n_459), .B(n_453), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_457), .B(n_432), .C(n_443), .Y(n_463) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_458), .A2(n_446), .B(n_447), .C(n_454), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_462), .B(n_455), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_463), .Y(n_466) );
XNOR2xp5_ASAP7_75t_L g467 ( .A(n_461), .B(n_456), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_466), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_467), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_469), .B(n_464), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_470), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_471), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_472), .A2(n_465), .B(n_468), .Y(n_473) );
endmodule