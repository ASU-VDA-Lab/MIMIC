module fake_jpeg_24444_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_38),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx11_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_27),
.B1(n_36),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_76),
.B1(n_80),
.B2(n_30),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_35),
.B(n_31),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_60),
.Y(n_101)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_69),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_78),
.Y(n_97)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_19),
.B1(n_22),
.B2(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_15),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_26),
.B1(n_32),
.B2(n_19),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_89),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_57),
.Y(n_120)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_35),
.B1(n_30),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_117),
.B1(n_80),
.B2(n_86),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_115),
.B1(n_79),
.B2(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_26),
.Y(n_127)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_56),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_20),
.B(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_130),
.B1(n_132),
.B2(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_73),
.Y(n_128)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_134),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_68),
.B1(n_56),
.B2(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_84),
.B1(n_77),
.B2(n_23),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_102),
.B1(n_105),
.B2(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_77),
.Y(n_135)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_13),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_13),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_1),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_93),
.B1(n_106),
.B2(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_1),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_2),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_104),
.C(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_133),
.B1(n_122),
.B2(n_129),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_162),
.Y(n_181)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_104),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_108),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_127),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_4),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_173),
.C(n_143),
.Y(n_187)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_5),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_11),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_138),
.B(n_147),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_176),
.B1(n_169),
.B2(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_161),
.A2(n_140),
.B(n_137),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_173),
.C(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_121),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_136),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_158),
.B(n_145),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_132),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_176),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_151),
.B(n_168),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_205),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_210),
.B1(n_186),
.B2(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_194),
.B1(n_190),
.B2(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_148),
.B1(n_90),
.B2(n_124),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_160),
.C(n_152),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_154),
.A3(n_171),
.B1(n_163),
.B2(n_156),
.C1(n_90),
.C2(n_124),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_222),
.B(n_223),
.C(n_225),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_191),
.B(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_199),
.B1(n_201),
.B2(n_200),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_227),
.A2(n_202),
.B1(n_179),
.B2(n_155),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_220),
.Y(n_245)
);

NAND4xp25_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_202),
.C(n_199),
.D(n_156),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_211),
.C(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_238),
.C(n_218),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_203),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_212),
.C(n_10),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_246),
.C(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_248),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_225),
.B1(n_222),
.B2(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_216),
.B1(n_229),
.B2(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_231),
.B(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_246),
.C(n_230),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_230),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_248),
.B(n_217),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_249),
.A2(n_241),
.B1(n_251),
.B2(n_252),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_5),
.B(n_6),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_5),
.B(n_6),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.C(n_260),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_255),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_264),
.B(n_7),
.CI(n_8),
.CON(n_265),
.SN(n_265)
);


endmodule