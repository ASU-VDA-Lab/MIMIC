module fake_netlist_6_803_n_111 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_111);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_111;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_85;
wire n_66;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp67_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_R g54 ( 
.A(n_53),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_34),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_42),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_37),
.Y(n_60)
);

OR2x6_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_25),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_R g64 ( 
.A(n_59),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_57),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_45),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_40),
.B(n_42),
.C(n_23),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_61),
.B1(n_37),
.B2(n_60),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_61),
.B1(n_38),
.B2(n_64),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_61),
.B1(n_68),
.B2(n_71),
.C(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_64),
.B1(n_69),
.B2(n_37),
.Y(n_78)
);

AO21x2_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_69),
.B(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_20),
.C(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_12),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_16),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_15),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_77),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_79),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_84),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_84),
.B(n_85),
.C(n_82),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_81),
.B1(n_85),
.B2(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_90),
.Y(n_96)
);

AOI211xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_94),
.B(n_21),
.C(n_34),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_3),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_R g100 ( 
.A(n_98),
.B(n_6),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_97),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_6),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_7),
.Y(n_103)
);

AOI222xp33_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_34),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_37),
.Y(n_104)
);

NAND4xp25_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_100),
.C(n_8),
.D(n_50),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

OAI211xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_34),
.B(n_37),
.C(n_52),
.Y(n_107)
);

NAND4xp75_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_106),
.C(n_52),
.D(n_50),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_60),
.A3(n_37),
.B1(n_51),
.B2(n_49),
.C1(n_48),
.C2(n_47),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_49),
.B1(n_51),
.B2(n_48),
.C(n_47),
.Y(n_111)
);


endmodule