module fake_jpeg_10946_n_636 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_636);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_636;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_63),
.B(n_71),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_67),
.Y(n_166)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_10),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_72),
.Y(n_160)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_29),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_16),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_120),
.Y(n_127)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_20),
.B(n_11),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_109),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_11),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_45),
.C(n_47),
.Y(n_182)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_122),
.C(n_123),
.Y(n_146)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_21),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_121),
.A2(n_54),
.B1(n_44),
.B2(n_42),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_44),
.B1(n_54),
.B2(n_21),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_58),
.B1(n_57),
.B2(n_28),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_58),
.B1(n_57),
.B2(n_56),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_58),
.B1(n_57),
.B2(n_56),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_20),
.B1(n_55),
.B2(n_40),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_139),
.A2(n_149),
.B1(n_177),
.B2(n_35),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_140),
.B(n_189),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_20),
.B1(n_55),
.B2(n_40),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_36),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_168),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_86),
.A2(n_53),
.B1(n_21),
.B2(n_50),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_163),
.A2(n_197),
.B1(n_34),
.B2(n_74),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_53),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_60),
.B(n_50),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_170),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_48),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_65),
.B(n_25),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_175),
.B(n_176),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_45),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_91),
.A2(n_55),
.B1(n_24),
.B2(n_47),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_89),
.B(n_48),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_192),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_16),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_42),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_109),
.B(n_42),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_90),
.B(n_24),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_199),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_92),
.A2(n_54),
.B1(n_44),
.B2(n_33),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_62),
.B(n_42),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_84),
.A2(n_42),
.B1(n_39),
.B2(n_33),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_84),
.B1(n_69),
.B2(n_88),
.Y(n_214)
);

CKINVDCx6p67_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_204),
.Y(n_297)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_94),
.B1(n_103),
.B2(n_96),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_207),
.A2(n_243),
.B1(n_273),
.B2(n_184),
.Y(n_281)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_208),
.Y(n_306)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_209),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_211),
.B(n_250),
.Y(n_305)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_212),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_214),
.A2(n_234),
.B1(n_237),
.B2(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_215),
.Y(n_323)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_216),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_125),
.A2(n_121),
.B1(n_112),
.B2(n_105),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_218),
.A2(n_222),
.B1(n_232),
.B2(n_166),
.Y(n_325)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_139),
.A2(n_101),
.B1(n_70),
.B2(n_95),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g294 ( 
.A1(n_220),
.A2(n_264),
.B1(n_143),
.B2(n_126),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_182),
.A2(n_100),
.B1(n_85),
.B2(n_39),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_221),
.A2(n_180),
.B(n_132),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_149),
.A2(n_68),
.B1(n_66),
.B2(n_64),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_254),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_117),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_225),
.B(n_248),
.Y(n_291)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_226),
.Y(n_335)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_144),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_134),
.A2(n_73),
.B1(n_67),
.B2(n_61),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_126),
.A2(n_116),
.B1(n_104),
.B2(n_13),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_147),
.Y(n_240)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_201),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

NAND2x1_ASAP7_75t_L g253 ( 
.A(n_136),
.B(n_104),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_35),
.Y(n_319)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_255),
.B(n_268),
.Y(n_298)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_256),
.B(n_257),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_177),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_260),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_153),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_133),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_263),
.Y(n_309)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_35),
.B1(n_9),
.B2(n_12),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_127),
.B(n_12),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_277),
.Y(n_279)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_142),
.A2(n_137),
.B(n_124),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_267),
.B(n_270),
.Y(n_326)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_146),
.A2(n_35),
.B(n_7),
.C(n_14),
.D(n_18),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_160),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_271),
.Y(n_307)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_272),
.B(n_274),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_141),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_153),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_202),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_14),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_281),
.A2(n_220),
.B1(n_274),
.B2(n_247),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_198),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_288),
.B(n_289),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_249),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_225),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_290),
.B(n_310),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_219),
.A2(n_186),
.B1(n_198),
.B2(n_184),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_292),
.A2(n_316),
.B1(n_325),
.B2(n_330),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_294),
.B(n_304),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_213),
.B(n_151),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_295),
.B(n_332),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_224),
.B(n_154),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_217),
.A2(n_151),
.A3(n_150),
.B1(n_155),
.B2(n_152),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_210),
.A2(n_186),
.B1(n_191),
.B2(n_135),
.Y(n_312)
);

AO21x2_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_273),
.B(n_204),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_267),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_204),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_210),
.A2(n_166),
.B1(n_155),
.B2(n_150),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_324),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_222),
.A2(n_171),
.B1(n_135),
.B2(n_202),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_223),
.B(n_171),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_218),
.A2(n_180),
.B1(n_152),
.B2(n_132),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_340),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_221),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_207),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_214),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_340)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_355),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_281),
.A2(n_220),
.B1(n_237),
.B2(n_234),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_345),
.A2(n_342),
.B1(n_351),
.B2(n_381),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_326),
.A2(n_208),
.B(n_215),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_346),
.A2(n_357),
.B(n_323),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_347),
.A2(n_379),
.B1(n_297),
.B2(n_334),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_291),
.A2(n_268),
.B(n_264),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_348),
.A2(n_369),
.B(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_289),
.B(n_254),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_377),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_326),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_351),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_326),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_279),
.B(n_264),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_353),
.B(n_362),
.Y(n_421)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_262),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_302),
.A2(n_275),
.B(n_259),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_358),
.Y(n_393)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_314),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_371),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_278),
.B1(n_339),
.B2(n_320),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_295),
.B(n_216),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_366),
.Y(n_409)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_367),
.B(n_374),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_304),
.B(n_250),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_368),
.B(n_386),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_209),
.B(n_244),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_288),
.B(n_246),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_309),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_321),
.A2(n_231),
.B(n_239),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_304),
.B(n_205),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_376),
.B(n_382),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_332),
.B(n_302),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_383),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_298),
.A2(n_266),
.B1(n_271),
.B2(n_238),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_292),
.A2(n_229),
.B1(n_15),
.B2(n_17),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_380),
.A2(n_308),
.B1(n_300),
.B2(n_313),
.Y(n_395)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_283),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_283),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_389),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_302),
.B(n_229),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_336),
.A2(n_260),
.B1(n_15),
.B2(n_4),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_388),
.A2(n_318),
.B1(n_323),
.B2(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_286),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_356),
.A2(n_310),
.B1(n_294),
.B2(n_324),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_373),
.A2(n_294),
.B1(n_330),
.B2(n_337),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_373),
.A2(n_294),
.B1(n_307),
.B2(n_329),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_384),
.B1(n_381),
.B2(n_379),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_294),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_400),
.A2(n_348),
.B(n_374),
.Y(n_446)
);

OA22x2_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_406),
.B1(n_380),
.B2(n_361),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_296),
.B1(n_286),
.B2(n_300),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_404),
.A2(n_412),
.B1(n_361),
.B2(n_402),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_306),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_428),
.B(n_399),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_349),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_417),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_305),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_422),
.C(n_425),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_360),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_296),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_342),
.A2(n_287),
.B(n_339),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_369),
.B(n_346),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_333),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_341),
.B(n_284),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_341),
.Y(n_438)
);

AOI21xp33_ASAP7_75t_SL g428 ( 
.A1(n_384),
.A2(n_287),
.B(n_306),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_344),
.B(n_284),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_429),
.B(n_411),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_386),
.C(n_378),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_433),
.B(n_443),
.C(n_451),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_435),
.A2(n_446),
.B(n_455),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_436),
.A2(n_445),
.B1(n_465),
.B2(n_404),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_420),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_440),
.Y(n_475)
);

OAI221xp5_ASAP7_75t_SL g495 ( 
.A1(n_438),
.A2(n_458),
.B1(n_460),
.B2(n_462),
.C(n_401),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_422),
.B(n_384),
.Y(n_439)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_413),
.B(n_383),
.Y(n_441)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_405),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_442),
.B(n_468),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_357),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_450),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_353),
.B1(n_361),
.B2(n_371),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_365),
.Y(n_447)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_448),
.B(n_429),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_449),
.A2(n_459),
.B1(n_466),
.B2(n_410),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_367),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_421),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_421),
.C(n_441),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_372),
.B(n_352),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_464),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_397),
.B(n_358),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_400),
.A2(n_361),
.B1(n_375),
.B2(n_382),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_389),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_430),
.A2(n_364),
.B1(n_354),
.B2(n_377),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_430),
.B1(n_428),
.B2(n_407),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_385),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_405),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_398),
.A2(n_361),
.B1(n_375),
.B2(n_364),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_400),
.A2(n_278),
.B1(n_343),
.B2(n_359),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_333),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_425),
.C(n_408),
.Y(n_476)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_469),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_471),
.B(n_472),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_448),
.B(n_432),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_474),
.B(n_501),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_478),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_477),
.A2(n_450),
.B1(n_418),
.B2(n_403),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_432),
.B(n_414),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_481),
.A2(n_484),
.B1(n_493),
.B2(n_430),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_434),
.A2(n_465),
.B1(n_445),
.B2(n_436),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_414),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_488),
.B(n_492),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_426),
.C(n_410),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_491),
.C(n_496),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_426),
.C(n_410),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_426),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_434),
.A2(n_442),
.B1(n_440),
.B2(n_437),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_444),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_495),
.B(n_499),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_446),
.C(n_438),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_408),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_500),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_454),
.A2(n_423),
.B(n_431),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_394),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_452),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_410),
.C(n_431),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_503),
.C(n_435),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_418),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_463),
.Y(n_504)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_505),
.B(n_522),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_482),
.A2(n_455),
.B1(n_458),
.B2(n_460),
.Y(n_507)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_466),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_509),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_510),
.A2(n_390),
.B1(n_317),
.B2(n_299),
.Y(n_548)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_511),
.A2(n_517),
.B1(n_523),
.B2(n_524),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_514),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_478),
.B(n_459),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_449),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_519),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_470),
.A2(n_469),
.B(n_468),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_516),
.A2(n_520),
.B(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_457),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_499),
.A2(n_470),
.B(n_489),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_456),
.B(n_450),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_415),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_493),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_528),
.A2(n_481),
.B1(n_484),
.B2(n_489),
.Y(n_537)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_529),
.B(n_479),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_403),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_280),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_471),
.B(n_395),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_532),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_472),
.B(n_450),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_533),
.A2(n_477),
.B1(n_502),
.B2(n_496),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_473),
.C(n_490),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_534),
.B(n_535),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_530),
.C(n_512),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_537),
.A2(n_328),
.B1(n_285),
.B2(n_335),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_538),
.A2(n_547),
.B1(n_554),
.B2(n_531),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_480),
.Y(n_541)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_541),
.Y(n_572)
);

CKINVDCx14_ASAP7_75t_R g570 ( 
.A(n_544),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_497),
.Y(n_546)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_546),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_533),
.A2(n_494),
.B1(n_473),
.B2(n_492),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_553),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_390),
.C(n_293),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_551),
.C(n_555),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_282),
.Y(n_550)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_550),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_513),
.B(n_293),
.C(n_282),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_526),
.A2(n_317),
.B1(n_280),
.B2(n_311),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_514),
.B(n_328),
.C(n_285),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_518),
.B(n_525),
.C(n_519),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_558),
.A2(n_520),
.B(n_526),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_559),
.A2(n_562),
.B(n_536),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_550),
.A2(n_521),
.B1(n_516),
.B2(n_504),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_566),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_547),
.A2(n_510),
.B1(n_528),
.B2(n_532),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_574),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_558),
.A2(n_510),
.B(n_525),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_557),
.B(n_518),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_564),
.B(n_556),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g587 ( 
.A(n_565),
.B(n_536),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_541),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_508),
.Y(n_567)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_567),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_508),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_568),
.B(n_572),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_569),
.A2(n_579),
.B1(n_549),
.B2(n_551),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_538),
.A2(n_260),
.B1(n_335),
.B2(n_15),
.Y(n_574)
);

BUFx24_ASAP7_75t_SL g577 ( 
.A(n_542),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_553),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_555),
.Y(n_579)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_559),
.A2(n_573),
.B(n_571),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_582),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_535),
.C(n_539),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_575),
.B(n_539),
.C(n_534),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_583),
.B(n_588),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_585),
.B(n_587),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_565),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_590),
.B(n_593),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_545),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_591),
.B(n_595),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_572),
.A2(n_554),
.B1(n_552),
.B2(n_537),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_594),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_573),
.A2(n_548),
.B1(n_545),
.B2(n_4),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_578),
.B(n_0),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_3),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_595),
.Y(n_600)
);

OAI211xp5_ASAP7_75t_SL g608 ( 
.A1(n_597),
.A2(n_568),
.B(n_576),
.C(n_579),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_600),
.B(n_596),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_570),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_610),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_582),
.B(n_576),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_606),
.B(n_609),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_561),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_607),
.B(n_584),
.C(n_4),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_6),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_583),
.B(n_562),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_569),
.C(n_574),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_589),
.C(n_586),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_612),
.B(n_615),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_603),
.A2(n_597),
.B(n_587),
.Y(n_613)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_613),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_614),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_611),
.A2(n_584),
.B(n_4),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_618),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_6),
.C(n_610),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_617),
.B(n_600),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_599),
.B(n_6),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_621),
.B(n_6),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_SL g628 ( 
.A1(n_625),
.A2(n_618),
.B(n_620),
.C(n_619),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_626),
.B(n_598),
.C(n_617),
.Y(n_630)
);

NAND2x1_ASAP7_75t_L g632 ( 
.A(n_628),
.B(n_627),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_622),
.A2(n_612),
.B(n_604),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_629),
.B(n_630),
.C(n_623),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_632),
.C(n_623),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_632),
.C(n_601),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_624),
.C(n_601),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_598),
.B(n_6),
.Y(n_636)
);


endmodule