module fake_jpeg_28895_n_446 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_446);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_8),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_48),
.B(n_52),
.Y(n_130)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_53),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g108 ( 
.A(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_64),
.Y(n_124)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_0),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_7),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_72),
.C(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_79),
.B(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_21),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_19),
.B1(n_20),
.B2(n_38),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_93),
.A2(n_55),
.B1(n_19),
.B2(n_82),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_22),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_104),
.B(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_51),
.Y(n_142)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_62),
.B(n_43),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_46),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_72),
.B(n_69),
.C(n_35),
.Y(n_139)
);

NOR2x1_ASAP7_75t_R g193 ( 
.A(n_139),
.B(n_30),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx2_ASAP7_75t_SL g200 ( 
.A(n_140),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_148),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_147),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_21),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_133),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_25),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_162),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_158),
.B1(n_67),
.B2(n_71),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_22),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_160),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_22),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_47),
.B1(n_63),
.B2(n_66),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_171),
.B1(n_172),
.B2(n_103),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_85),
.B1(n_77),
.B2(n_78),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_51),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_25),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_111),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_30),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_105),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_100),
.B(n_115),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_123),
.B(n_94),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_88),
.B1(n_114),
.B2(n_119),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_190),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_108),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_155),
.C(n_136),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_94),
.B(n_110),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_110),
.B(n_95),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_105),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_196),
.B1(n_96),
.B2(n_91),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_R g214 ( 
.A(n_193),
.B(n_157),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_119),
.B1(n_106),
.B2(n_109),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_204),
.B(n_211),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_205),
.A2(n_189),
.B(n_180),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_208),
.B1(n_163),
.B2(n_151),
.Y(n_244)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_192),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_143),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_178),
.B(n_30),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_221),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_225),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_109),
.B1(n_141),
.B2(n_68),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_184),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_74),
.B1(n_54),
.B2(n_56),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_61),
.B1(n_96),
.B2(n_118),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_169),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_175),
.B(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_153),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_152),
.C(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_199),
.C(n_192),
.Y(n_231)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_224),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_165),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_236),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_234),
.B(n_246),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_188),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_235),
.C(n_250),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_202),
.C(n_199),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_179),
.C(n_173),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_186),
.B1(n_197),
.B2(n_181),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_91),
.B1(n_90),
.B2(n_118),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_200),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_227),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_210),
.B(n_176),
.CI(n_197),
.CON(n_249),
.SN(n_249)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_226),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_206),
.A2(n_214),
.B1(n_205),
.B2(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_253),
.A2(n_146),
.B1(n_137),
.B2(n_102),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

CKINVDCx12_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_257),
.A2(n_259),
.B(n_265),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_263),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_223),
.C(n_207),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_231),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_227),
.B(n_208),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_273),
.Y(n_295)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_217),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_227),
.B(n_216),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_278),
.B(n_177),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_230),
.B(n_238),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_159),
.B(n_220),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_279),
.A2(n_195),
.B1(n_198),
.B2(n_194),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_251),
.B1(n_241),
.B2(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_282),
.A2(n_286),
.B1(n_298),
.B2(n_274),
.Y(n_327)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_236),
.B1(n_245),
.B2(n_249),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_285),
.A2(n_303),
.B(n_252),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_240),
.B1(n_229),
.B2(n_230),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_249),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_253),
.B(n_235),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_291),
.B(n_263),
.CI(n_171),
.CON(n_330),
.SN(n_330)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_261),
.C(n_264),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_258),
.B(n_220),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_301),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_195),
.B1(n_194),
.B2(n_198),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_272),
.B1(n_278),
.B2(n_262),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_254),
.B(n_12),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_306),
.B(n_265),
.Y(n_311)
);

AO22x1_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_198),
.B1(n_144),
.B2(n_164),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_277),
.B(n_266),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_260),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_177),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_255),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_257),
.A2(n_149),
.B(n_146),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_272),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_252),
.A2(n_33),
.B1(n_38),
.B2(n_90),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_261),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_330),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.C(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_264),
.C(n_255),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_273),
.B1(n_271),
.B2(n_259),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_329),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_303),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_285),
.A2(n_271),
.B(n_276),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_295),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_268),
.B1(n_267),
.B2(n_279),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_263),
.C(n_137),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_0),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_332),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_300),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_161),
.C(n_131),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.C(n_298),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_131),
.C(n_126),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_286),
.C(n_306),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_339),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_346),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_307),
.B1(n_308),
.B2(n_285),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_282),
.C(n_280),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_347),
.C(n_348),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_287),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_287),
.C(n_295),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_290),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_284),
.B1(n_292),
.B2(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_11),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_302),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_357),
.C(n_331),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_356),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_288),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_288),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_332),
.B(n_38),
.CI(n_33),
.CON(n_358),
.SN(n_358)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_318),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_344),
.A2(n_319),
.B(n_322),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_317),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_368),
.Y(n_382)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_330),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_367),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_316),
.C(n_322),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_357),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_375),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_376),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_354),
.A2(n_323),
.B(n_333),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_373),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_353),
.A2(n_334),
.B1(n_126),
.B2(n_106),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_41),
.Y(n_375)
);

AO221x1_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_35),
.B1(n_171),
.B2(n_13),
.C(n_18),
.Y(n_376)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_377),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_SL g383 ( 
.A1(n_378),
.A2(n_379),
.B(n_17),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_12),
.B(n_18),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_335),
.C(n_341),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_385),
.Y(n_399)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_375),
.A2(n_352),
.B1(n_338),
.B2(n_340),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_372),
.C(n_359),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_335),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_388),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_10),
.B1(n_17),
.B2(n_12),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_33),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_379),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_360),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_382),
.B(n_362),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_397),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_372),
.C(n_391),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_401),
.C(n_375),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_370),
.C(n_371),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_390),
.B(n_367),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_172),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_393),
.A2(n_361),
.B(n_367),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_407),
.A2(n_395),
.B(n_390),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_392),
.B(n_365),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_377),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_412),
.Y(n_428)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_399),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_411),
.B(n_420),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_378),
.C(n_395),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_402),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_414),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_383),
.C(n_76),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_415),
.A2(n_418),
.B(n_406),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_9),
.B(n_17),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_406),
.B(n_1),
.Y(n_423)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_84),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_405),
.A2(n_105),
.B(n_84),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_9),
.Y(n_420)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_423),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_417),
.C(n_76),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_0),
.B(n_1),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_426),
.A2(n_427),
.B(n_2),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_1),
.B(n_2),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_415),
.B(n_2),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_3),
.B(n_4),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_424),
.C(n_27),
.Y(n_438)
);

AOI322xp5_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_5),
.A3(n_6),
.B1(n_27),
.B2(n_377),
.C1(n_398),
.C2(n_364),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_425),
.C(n_429),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_434),
.A2(n_3),
.B(n_5),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_438),
.Y(n_441)
);

XOR2x2_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_440),
.Y(n_442)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_436),
.B(n_431),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_441),
.Y(n_444)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_444),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_6),
.Y(n_446)
);


endmodule