module real_aes_2352_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_171;
wire n_87;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_0), .A2(n_75), .B1(n_146), .B2(n_149), .Y(n_145) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_1), .A2(n_53), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g197 ( .A(n_2), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_3), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g254 ( .A(n_4), .Y(n_254) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_5), .A2(n_20), .B1(n_91), .B2(n_95), .Y(n_94) );
AOI22xp5_ASAP7_75t_L g85 ( .A1(n_6), .A2(n_8), .B1(n_86), .B2(n_104), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_7), .Y(n_269) );
INVx2_ASAP7_75t_L g217 ( .A(n_9), .Y(n_217) );
INVx1_ASAP7_75t_L g288 ( .A(n_10), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_11), .A2(n_49), .B1(n_124), .B2(n_132), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_12), .A2(n_72), .B1(n_111), .B2(n_118), .Y(n_110) );
INVx1_ASAP7_75t_L g285 ( .A(n_13), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_14), .A2(n_81), .B1(n_82), .B2(n_170), .Y(n_80) );
INVx1_ASAP7_75t_L g170 ( .A(n_14), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_15), .A2(n_47), .B1(n_136), .B2(n_140), .Y(n_135) );
INVx1_ASAP7_75t_SL g339 ( .A(n_16), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_17), .B(n_237), .Y(n_301) );
AOI33xp33_ASAP7_75t_L g325 ( .A1(n_18), .A2(n_38), .A3(n_222), .B1(n_230), .B2(n_326), .B3(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g262 ( .A(n_19), .Y(n_262) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_20), .A2(n_53), .B1(n_57), .B2(n_190), .C(n_192), .Y(n_189) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_21), .A2(n_68), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g247 ( .A(n_21), .B(n_68), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_22), .B(n_220), .Y(n_336) );
INVx3_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
AOI222xp33_ASAP7_75t_L g158 ( .A1(n_24), .A2(n_56), .B1(n_65), .B2(n_159), .C1(n_162), .C2(n_167), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_25), .A2(n_69), .B1(n_175), .B2(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_25), .Y(n_176) );
INVx1_ASAP7_75t_SL g99 ( .A(n_26), .Y(n_99) );
INVx1_ASAP7_75t_L g199 ( .A(n_27), .Y(n_199) );
AND2x2_ASAP7_75t_L g225 ( .A(n_27), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g243 ( .A(n_27), .B(n_197), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_28), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_29), .B(n_220), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_30), .A2(n_215), .B1(n_279), .B2(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_31), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_32), .B(n_237), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_33), .B(n_251), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_34), .B(n_237), .Y(n_255) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_35), .A2(n_57), .B1(n_91), .B2(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_36), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_37), .A2(n_173), .B1(n_174), .B2(n_177), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_37), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_39), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g223 ( .A(n_40), .Y(n_223) );
INVx1_ASAP7_75t_L g239 ( .A(n_40), .Y(n_239) );
AND2x2_ASAP7_75t_L g244 ( .A(n_41), .B(n_245), .Y(n_244) );
XOR2xp5_ASAP7_75t_L g584 ( .A(n_42), .B(n_81), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_43), .A2(n_59), .B1(n_220), .B2(n_228), .C(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_44), .B(n_220), .Y(n_313) );
INVx1_ASAP7_75t_L g100 ( .A(n_45), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_46), .B(n_215), .Y(n_271) );
AOI21xp5_ASAP7_75t_SL g309 ( .A1(n_48), .A2(n_228), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g282 ( .A(n_50), .Y(n_282) );
INVx1_ASAP7_75t_L g234 ( .A(n_51), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_52), .A2(n_228), .B(n_233), .Y(n_227) );
INVxp33_ASAP7_75t_L g194 ( .A(n_53), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_54), .A2(n_73), .B1(n_153), .B2(n_156), .Y(n_152) );
INVx1_ASAP7_75t_L g226 ( .A(n_55), .Y(n_226) );
INVx1_ASAP7_75t_L g241 ( .A(n_55), .Y(n_241) );
INVxp67_ASAP7_75t_L g193 ( .A(n_57), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_58), .B(n_220), .Y(n_328) );
INVx1_ASAP7_75t_L g183 ( .A(n_59), .Y(n_183) );
AND2x2_ASAP7_75t_L g341 ( .A(n_60), .B(n_214), .Y(n_341) );
INVx1_ASAP7_75t_L g283 ( .A(n_61), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_62), .A2(n_228), .B(n_338), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_62), .A2(n_81), .B1(n_82), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_62), .Y(n_577) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_63), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_63), .A2(n_228), .B(n_300), .C(n_304), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_64), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_64), .Y(n_179) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_66), .B(n_214), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_67), .A2(n_228), .B1(n_323), .B2(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g175 ( .A(n_69), .Y(n_175) );
INVx1_ASAP7_75t_L g311 ( .A(n_70), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_71), .B(n_214), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_74), .A2(n_260), .B(n_261), .C(n_264), .Y(n_259) );
BUFx2_ASAP7_75t_SL g191 ( .A(n_76), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_77), .B(n_237), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_186), .B1(n_200), .B2(n_571), .C(n_575), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_171), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND4xp75_ASAP7_75t_L g83 ( .A(n_84), .B(n_122), .C(n_144), .D(n_158), .Y(n_83) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_110), .Y(n_84) );
INVx4_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
AND2x2_ASAP7_75t_L g139 ( .A(n_89), .B(n_116), .Y(n_139) );
AND2x4_ASAP7_75t_L g151 ( .A(n_89), .B(n_131), .Y(n_151) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
INVx2_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
AND2x2_ASAP7_75t_L g143 ( .A(n_90), .B(n_94), .Y(n_143) );
INVx1_ASAP7_75t_L g92 ( .A(n_91), .Y(n_92) );
INVx2_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
OAI22x1_ASAP7_75t_L g97 ( .A1(n_91), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_91), .Y(n_98) );
INVx1_ASAP7_75t_L g103 ( .A(n_91), .Y(n_103) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x4_ASAP7_75t_L g114 ( .A(n_94), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
AND2x4_ASAP7_75t_L g155 ( .A(n_96), .B(n_129), .Y(n_155) );
AND2x2_ASAP7_75t_L g161 ( .A(n_96), .B(n_114), .Y(n_161) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_101), .Y(n_96) );
AND2x2_ASAP7_75t_L g107 ( .A(n_97), .B(n_102), .Y(n_107) );
INVx2_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_97), .Y(n_166) );
AND2x4_ASAP7_75t_L g131 ( .A(n_101), .B(n_117), .Y(n_131) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g116 ( .A(n_102), .B(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
BUFx6f_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x4_ASAP7_75t_L g120 ( .A(n_107), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g169 ( .A(n_107), .B(n_129), .Y(n_169) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
AND2x4_ASAP7_75t_L g134 ( .A(n_114), .B(n_131), .Y(n_134) );
INVxp67_ASAP7_75t_L g121 ( .A(n_115), .Y(n_121) );
AND2x4_ASAP7_75t_L g129 ( .A(n_115), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g148 ( .A(n_116), .B(n_129), .Y(n_148) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx6_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_135), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
AND2x4_ASAP7_75t_L g157 ( .A(n_131), .B(n_143), .Y(n_157) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g165 ( .A(n_143), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_152), .Y(n_144) );
INVx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx6_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
XNOR2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_178), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_174), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_184), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
AND3x1_ASAP7_75t_SL g188 ( .A(n_189), .B(n_195), .C(n_198), .Y(n_188) );
INVxp67_ASAP7_75t_L g583 ( .A(n_189), .Y(n_583) );
CKINVDCx8_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_195), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_195), .A2(n_296), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g221 ( .A(n_196), .B(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_SL g587 ( .A(n_196), .B(n_198), .Y(n_587) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g232 ( .A(n_197), .B(n_223), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_198), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g229 ( .A(n_199), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND4xp75_ASAP7_75t_L g203 ( .A(n_204), .B(n_443), .C(n_488), .D(n_557), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_403), .Y(n_205) );
NOR3xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_359), .C(n_384), .Y(n_206) );
OAI222xp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_273), .B1(n_314), .B2(n_330), .C1(n_346), .C2(n_353), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_248), .Y(n_209) );
AND2x2_ASAP7_75t_L g568 ( .A(n_210), .B(n_382), .Y(n_568) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_212), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_212), .B(n_257), .Y(n_358) );
INVx3_ASAP7_75t_L g373 ( .A(n_212), .Y(n_373) );
AND2x2_ASAP7_75t_L g506 ( .A(n_212), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_218), .B(n_244), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_214), .B1(n_259), .B2(n_265), .Y(n_258) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_213), .A2(n_218), .B(n_244), .Y(n_391) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_215), .B(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx4f_ASAP7_75t_L g251 ( .A(n_216), .Y(n_251) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_217), .B(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g279 ( .A(n_217), .B(n_247), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
INVx1_ASAP7_75t_L g272 ( .A(n_220), .Y(n_272) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_224), .Y(n_220) );
INVx1_ASAP7_75t_L g296 ( .A(n_221), .Y(n_296) );
OR2x6_ASAP7_75t_L g235 ( .A(n_222), .B(n_231), .Y(n_235) );
INVxp33_ASAP7_75t_L g326 ( .A(n_222), .Y(n_326) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g290 ( .A(n_223), .B(n_240), .Y(n_290) );
INVx1_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
BUFx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x6_ASAP7_75t_L g574 ( .A(n_225), .B(n_232), .Y(n_574) );
INVx2_ASAP7_75t_L g231 ( .A(n_226), .Y(n_231) );
AND2x6_ASAP7_75t_L g287 ( .A(n_226), .B(n_238), .Y(n_287) );
INVxp67_ASAP7_75t_L g270 ( .A(n_228), .Y(n_270) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_232), .Y(n_228) );
INVx1_ASAP7_75t_L g327 ( .A(n_230), .Y(n_327) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_242), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_235), .A2(n_242), .B(n_254), .C(n_255), .Y(n_253) );
INVxp67_ASAP7_75t_L g260 ( .A(n_235), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_235), .A2(n_263), .B1(n_282), .B2(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g303 ( .A(n_235), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_235), .A2(n_242), .B(n_311), .C(n_312), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_SL g338 ( .A1(n_235), .A2(n_242), .B(n_339), .C(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g263 ( .A(n_237), .Y(n_263) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_242), .B(n_279), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_242), .A2(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g323 ( .A(n_242), .Y(n_323) );
INVx5_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_243), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_245), .Y(n_334) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g436 ( .A(n_248), .B(n_389), .Y(n_436) );
AND2x2_ASAP7_75t_L g438 ( .A(n_248), .B(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g473 ( .A(n_248), .Y(n_473) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_257), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_L g356 ( .A(n_250), .Y(n_356) );
INVx1_ASAP7_75t_L g375 ( .A(n_250), .Y(n_375) );
AND2x4_ASAP7_75t_L g382 ( .A(n_250), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_250), .B(n_320), .Y(n_398) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_250), .Y(n_507) );
INVx1_ASAP7_75t_L g517 ( .A(n_250), .Y(n_517) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_256), .Y(n_250) );
INVx2_ASAP7_75t_SL g304 ( .A(n_251), .Y(n_304) );
INVx1_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
INVx2_ASAP7_75t_L g370 ( .A(n_257), .Y(n_370) );
INVx1_ASAP7_75t_L g451 ( .A(n_257), .Y(n_451) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_266), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B1(n_271), .B2(n_272), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_275), .B(n_305), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_275), .B(n_332), .Y(n_426) );
INVx2_ASAP7_75t_L g447 ( .A(n_275), .Y(n_447) );
AND2x2_ASAP7_75t_L g455 ( .A(n_275), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_292), .Y(n_275) );
AND2x4_ASAP7_75t_L g345 ( .A(n_276), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g352 ( .A(n_276), .Y(n_352) );
AND2x2_ASAP7_75t_L g528 ( .A(n_276), .B(n_333), .Y(n_528) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g366 ( .A(n_277), .B(n_293), .Y(n_366) );
INVx2_ASAP7_75t_L g402 ( .A(n_277), .Y(n_402) );
AND2x2_ASAP7_75t_L g481 ( .A(n_277), .B(n_333), .Y(n_481) );
NOR2x1_ASAP7_75t_SL g524 ( .A(n_277), .B(n_306), .Y(n_524) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_279), .A2(n_309), .B(n_313), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B(n_291), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B1(n_288), .B2(n_289), .Y(n_284) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g364 ( .A(n_292), .Y(n_364) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g378 ( .A(n_293), .B(n_306), .Y(n_378) );
INVx1_ASAP7_75t_L g394 ( .A(n_293), .Y(n_394) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_293), .Y(n_502) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .C(n_298), .Y(n_295) );
INVxp67_ASAP7_75t_L g590 ( .A(n_297), .Y(n_590) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_304), .A2(n_321), .B(n_329), .Y(n_320) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_304), .A2(n_321), .B(n_329), .Y(n_371) );
AND2x2_ASAP7_75t_L g365 ( .A(n_305), .B(n_366), .Y(n_365) );
OR2x6_ASAP7_75t_L g446 ( .A(n_305), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g484 ( .A(n_305), .B(n_481), .Y(n_484) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx4_ASAP7_75t_L g343 ( .A(n_306), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_306), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g413 ( .A(n_306), .Y(n_413) );
OR2x2_ASAP7_75t_L g419 ( .A(n_306), .B(n_333), .Y(n_419) );
AND2x4_ASAP7_75t_L g433 ( .A(n_306), .B(n_394), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_306), .B(n_402), .Y(n_434) );
OR2x6_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g478 ( .A(n_317), .B(n_397), .Y(n_478) );
BUFx2_ASAP7_75t_L g530 ( .A(n_317), .Y(n_530) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g561 ( .A(n_319), .B(n_473), .Y(n_561) );
INVx2_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_328), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_342), .Y(n_330) );
AND2x2_ASAP7_75t_L g377 ( .A(n_331), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_SL g362 ( .A(n_332), .B(n_352), .Y(n_362) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g350 ( .A(n_333), .Y(n_350) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_333), .Y(n_456) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_333), .Y(n_523) );
INVx1_ASAP7_75t_L g563 ( .A(n_333), .Y(n_563) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B(n_341), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
OAI222xp33_ASAP7_75t_L g575 ( .A1(n_339), .A2(n_576), .B1(n_578), .B2(n_584), .C1(n_585), .C2(n_588), .Y(n_575) );
BUFx2_ASAP7_75t_L g477 ( .A(n_342), .Y(n_477) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x4_ASAP7_75t_L g393 ( .A(n_343), .B(n_394), .Y(n_393) );
NOR2xp67_ASAP7_75t_SL g425 ( .A(n_343), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g498 ( .A(n_343), .B(n_481), .Y(n_498) );
AND2x4_ASAP7_75t_SL g501 ( .A(n_343), .B(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g550 ( .A(n_343), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_345), .B(n_410), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_345), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_345), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g495 ( .A(n_349), .B(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g411 ( .A(n_350), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
AND2x2_ASAP7_75t_L g529 ( .A(n_354), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g537 ( .A(n_354), .B(n_466), .Y(n_537) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g406 ( .A(n_355), .B(n_391), .Y(n_406) );
AND2x4_ASAP7_75t_L g439 ( .A(n_355), .B(n_373), .Y(n_439) );
INVx1_ASAP7_75t_L g556 ( .A(n_355), .Y(n_556) );
AND2x2_ASAP7_75t_L g442 ( .A(n_357), .B(n_382), .Y(n_442) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g463 ( .A(n_358), .B(n_398), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_367), .B1(n_376), .B2(n_379), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_365), .Y(n_360) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_361), .A2(n_430), .B1(n_538), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_362), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g431 ( .A(n_362), .B(n_363), .Y(n_431) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_362), .B(n_433), .Y(n_461) );
AOI211xp5_ASAP7_75t_SL g549 ( .A1(n_362), .A2(n_550), .B(n_552), .C(n_553), .Y(n_549) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_363), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_363), .B(n_409), .Y(n_535) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g440 ( .A(n_365), .Y(n_440) );
INVx2_ASAP7_75t_L g496 ( .A(n_366), .Y(n_496) );
AND2x2_ASAP7_75t_L g570 ( .A(n_366), .B(n_563), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_367), .A2(n_519), .B(n_525), .Y(n_518) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g505 ( .A(n_369), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g515 ( .A(n_369), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g422 ( .A(n_370), .B(n_375), .Y(n_422) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_370), .B(n_391), .Y(n_424) );
AND2x2_ASAP7_75t_L g466 ( .A(n_370), .B(n_391), .Y(n_466) );
INVx2_ASAP7_75t_L g383 ( .A(n_371), .Y(n_383) );
AND2x4_ASAP7_75t_L g389 ( .A(n_371), .B(n_390), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx3_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
INVx3_ASAP7_75t_L g387 ( .A(n_374), .Y(n_387) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_378), .A2(n_484), .B(n_560), .Y(n_564) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g396 ( .A(n_381), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_381), .B(n_456), .Y(n_471) );
OR2x2_ASAP7_75t_L g486 ( .A(n_381), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g493 ( .A(n_381), .B(n_397), .Y(n_493) );
AND2x2_ASAP7_75t_L g449 ( .A(n_382), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g465 ( .A(n_382), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g482 ( .A(n_382), .B(n_451), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_392), .B1(n_395), .B2(n_399), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_387), .B(n_388), .Y(n_459) );
NOR2xp67_ASAP7_75t_SL g497 ( .A(n_387), .B(n_405), .Y(n_497) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_391), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g400 ( .A(n_393), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g464 ( .A(n_393), .B(n_410), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_393), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g567 ( .A(n_401), .B(n_433), .Y(n_567) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_402), .B(n_513), .Y(n_512) );
NOR2xp67_ASAP7_75t_SL g403 ( .A(n_404), .B(n_427), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B(n_414), .C(n_423), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_405), .A2(n_458), .B(n_468), .C(n_472), .Y(n_467) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g547 ( .A(n_406), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g458 ( .A(n_410), .B(n_434), .Y(n_458) );
AND2x2_ASAP7_75t_L g545 ( .A(n_410), .B(n_524), .Y(n_545) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g513 ( .A(n_413), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_420), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_417), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_435), .B1(n_437), .B2(n_440), .C(n_441), .Y(n_427) );
NOR4xp25_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .C(n_432), .D(n_434), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g546 ( .A(n_433), .B(n_509), .Y(n_546) );
INVx2_ASAP7_75t_L g552 ( .A(n_433), .Y(n_552) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_436), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g539 ( .A(n_439), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND4xp75_ASAP7_75t_L g444 ( .A(n_445), .B(n_467), .C(n_474), .D(n_483), .Y(n_444) );
OA211x2_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_452), .C(n_460), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_446), .B(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g540 ( .A(n_450), .Y(n_540) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g548 ( .A(n_451), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_459), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_464), .B2(n_465), .Y(n_460) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_464), .A2(n_515), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g543 ( .A(n_465), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_466), .B(n_556), .Y(n_555) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVxp67_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
AND2x2_ASAP7_75t_SL g500 ( .A(n_481), .B(n_501), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_482), .A2(n_545), .B1(n_567), .B2(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND3x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_531), .C(n_544), .Y(n_489) );
NOR3x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_503), .C(n_518), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_499), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_497), .B2(n_498), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_508), .B1(n_510), .B2(n_514), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g562 ( .A(n_512), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g551 ( .A(n_528), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_529), .A2(n_560), .B(n_562), .Y(n_559) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .B1(n_538), .B2(n_541), .Y(n_532) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
O2A1O1Ixp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_547), .C(n_549), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2x1_ASAP7_75t_SL g557 ( .A(n_558), .B(n_565), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .Y(n_558) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_566), .B(n_569), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
CKINVDCx16_ASAP7_75t_R g588 ( .A(n_589), .Y(n_588) );
endmodule