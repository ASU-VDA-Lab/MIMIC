module fake_jpeg_2176_n_504 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_504);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_504;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_51),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_1),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_53),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_57),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_62),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_2),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g155 ( 
.A(n_64),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_15),
.B(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_72),
.Y(n_107)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_69),
.B(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_14),
.B(n_5),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_85),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_96),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_25),
.A2(n_5),
.B(n_6),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_33),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_44),
.Y(n_137)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_151),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_44),
.B1(n_18),
.B2(n_29),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_106),
.A2(n_125),
.B1(n_140),
.B2(n_68),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_49),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_112),
.B1(n_118),
.B2(n_131),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_35),
.B1(n_24),
.B2(n_38),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_35),
.B1(n_46),
.B2(n_42),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g197 ( 
.A1(n_114),
.A2(n_126),
.B1(n_144),
.B2(n_145),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_44),
.B1(n_29),
.B2(n_31),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_53),
.A2(n_46),
.B1(n_42),
.B2(n_29),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_38),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_33),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_36),
.B1(n_39),
.B2(n_34),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_31),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_31),
.B1(n_29),
.B2(n_36),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_70),
.B(n_31),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_54),
.A2(n_39),
.B1(n_34),
.B2(n_26),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_40),
.B1(n_7),
.B2(n_8),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_29),
.Y(n_171)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_162),
.Y(n_225)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_163),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_109),
.A2(n_65),
.B1(n_59),
.B2(n_94),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_185),
.B1(n_140),
.B2(n_155),
.Y(n_219)
);

INVx5_ASAP7_75t_SL g166 ( 
.A(n_101),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_168),
.Y(n_241)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_171),
.B(n_173),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

AO22x2_ASAP7_75t_SL g177 ( 
.A1(n_114),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_177),
.A2(n_155),
.B(n_144),
.C(n_146),
.Y(n_236)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_78),
.B1(n_95),
.B2(n_93),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_180),
.A2(n_190),
.B1(n_191),
.B2(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_64),
.B1(n_88),
.B2(n_60),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_105),
.B(n_81),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_147),
.Y(n_212)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_139),
.A2(n_56),
.B1(n_63),
.B2(n_66),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_110),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_82),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_194),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_106),
.A2(n_89),
.B1(n_87),
.B2(n_83),
.Y(n_195)
);

AOI22x1_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_198),
.B1(n_200),
.B2(n_186),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_137),
.B(n_98),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_201),
.C(n_125),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_206),
.B1(n_131),
.B2(n_155),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g198 ( 
.A1(n_115),
.A2(n_71),
.B1(n_19),
.B2(n_79),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_108),
.A2(n_73),
.B1(n_19),
.B2(n_48),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_107),
.B(n_40),
.C(n_52),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_207),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_111),
.B(n_6),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_196),
.Y(n_224)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_197),
.B1(n_181),
.B2(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_208),
.A2(n_215),
.B1(n_240),
.B2(n_160),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_222),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_229),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_102),
.B1(n_103),
.B2(n_162),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_116),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_143),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_152),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_120),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_200),
.B(n_195),
.C(n_177),
.Y(n_246)
);

AND2x4_ASAP7_75t_SL g239 ( 
.A(n_196),
.B(n_157),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_143),
.B(n_157),
.C(n_102),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_113),
.B1(n_158),
.B2(n_146),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_197),
.B1(n_180),
.B2(n_177),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_248),
.B1(n_250),
.B2(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_195),
.B1(n_170),
.B2(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_198),
.B(n_170),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_268),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_113),
.B1(n_158),
.B2(n_145),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_263),
.B1(n_230),
.B2(n_219),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_176),
.B(n_166),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_179),
.B1(n_149),
.B2(n_127),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_149),
.B1(n_127),
.B2(n_150),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_266),
.B1(n_211),
.B2(n_225),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_178),
.B1(n_175),
.B2(n_163),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_205),
.B(n_202),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_270),
.B1(n_273),
.B2(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_123),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_271),
.Y(n_275)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_164),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_215),
.B1(n_232),
.B2(n_229),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_282),
.B1(n_283),
.B2(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_265),
.B1(n_247),
.B2(n_259),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_224),
.C(n_238),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_253),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_238),
.C(n_231),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_300),
.C(n_280),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_240),
.B1(n_231),
.B2(n_239),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_239),
.B1(n_236),
.B2(n_212),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_252),
.B(n_227),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_286),
.B(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_236),
.B1(n_227),
.B2(n_238),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_254),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_250),
.A2(n_211),
.B1(n_223),
.B2(n_199),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_262),
.A2(n_228),
.B1(n_223),
.B2(n_235),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_253),
.A2(n_223),
.B1(n_210),
.B2(n_234),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_256),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_249),
.A2(n_210),
.B1(n_243),
.B2(n_234),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_276),
.B1(n_289),
.B2(n_277),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_300),
.B(n_303),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_255),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_218),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_317),
.C(n_319),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_308),
.A2(n_322),
.B1(n_323),
.B2(n_326),
.Y(n_340)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_311),
.A2(n_320),
.B1(n_325),
.B2(n_225),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_267),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_318),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_316),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_271),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_269),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_269),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_285),
.A2(n_263),
.B1(n_244),
.B2(n_246),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_266),
.B1(n_264),
.B2(n_246),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_277),
.A2(n_269),
.B1(n_260),
.B2(n_261),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_265),
.B(n_245),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_265),
.B1(n_270),
.B2(n_268),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_274),
.A2(n_265),
.B(n_241),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_291),
.B1(n_283),
.B2(n_299),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_331),
.A2(n_278),
.B1(n_298),
.B2(n_287),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_273),
.B(n_225),
.Y(n_333)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_304),
.B(n_288),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_278),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_334),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_218),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_221),
.C(n_242),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_290),
.B1(n_279),
.B2(n_296),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_337),
.A2(n_342),
.B1(n_344),
.B2(n_348),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_275),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_349),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_332),
.A2(n_302),
.B1(n_301),
.B2(n_294),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_345),
.B1(n_350),
.B2(n_361),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_292),
.B1(n_304),
.B2(n_298),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_304),
.B1(n_292),
.B2(n_287),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_322),
.A2(n_273),
.B1(n_221),
.B2(n_242),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_213),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_358),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_314),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_327),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_213),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_209),
.B1(n_168),
.B2(n_190),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_331),
.A2(n_307),
.B1(n_326),
.B2(n_315),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_133),
.B1(n_123),
.B2(n_173),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_309),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_318),
.C(n_319),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.C(n_328),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_209),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_321),
.Y(n_368)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_355),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_335),
.C(n_328),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_382),
.C(n_384),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_340),
.A2(n_330),
.B1(n_307),
.B2(n_311),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_387),
.B1(n_361),
.B2(n_348),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_356),
.A2(n_333),
.B(n_321),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_383),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_328),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_377),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_316),
.Y(n_377)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_334),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_380),
.B(n_385),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_325),
.C(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_138),
.C(n_133),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_392),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_SL g388 ( 
.A(n_337),
.B(n_364),
.C(n_340),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_388),
.B(n_362),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_173),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_389),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_349),
.C(n_359),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_391),
.C(n_354),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_103),
.C(n_40),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_40),
.B(n_7),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_6),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_395),
.A2(n_400),
.B1(n_403),
.B2(n_375),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_401),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_353),
.B1(n_352),
.B2(n_336),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_408),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_393),
.A2(n_353),
.B1(n_352),
.B2(n_355),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_343),
.C(n_344),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_404),
.B(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_345),
.C(n_341),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_341),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_341),
.C(n_350),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_410),
.B(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_366),
.C(n_360),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_40),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_391),
.Y(n_437)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_415)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_6),
.C(n_8),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_378),
.C(n_389),
.Y(n_426)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_418),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_407),
.A2(n_368),
.B1(n_369),
.B2(n_374),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_SL g420 ( 
.A(n_412),
.B(n_367),
.C(n_389),
.Y(n_420)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_438),
.Y(n_441)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_429),
.Y(n_445)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_381),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_432),
.B(n_436),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_414),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_388),
.C(n_382),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_433),
.B(n_434),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_369),
.B1(n_387),
.B2(n_394),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_390),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_413),
.Y(n_452)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_398),
.C(n_404),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_444),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_424),
.A2(n_400),
.B1(n_405),
.B2(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_435),
.B(n_398),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_447),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_397),
.C(n_399),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_408),
.Y(n_448)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_397),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_451),
.B(n_453),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_8),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_417),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_14),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_8),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_421),
.A2(n_14),
.B1(n_9),
.B2(n_10),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_456),
.A2(n_422),
.B1(n_426),
.B2(n_437),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_425),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_457),
.B(n_468),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_429),
.A3(n_427),
.B1(n_421),
.B2(n_419),
.C(n_422),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_458),
.A2(n_455),
.B(n_452),
.Y(n_477)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_443),
.C(n_439),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_461),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_433),
.C(n_9),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_466),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_14),
.Y(n_478)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_449),
.B(n_10),
.CI(n_11),
.CON(n_466),
.SN(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_11),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_11),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_470),
.B(n_471),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_11),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_SL g472 ( 
.A(n_469),
.B(n_445),
.C(n_455),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_472),
.A2(n_473),
.B(n_466),
.C(n_468),
.Y(n_489)
);

AOI21x1_ASAP7_75t_L g473 ( 
.A1(n_464),
.A2(n_442),
.B(n_450),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_462),
.A2(n_442),
.B(n_445),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_477),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_481),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_12),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_12),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_13),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_461),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_486),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_457),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_490),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_480),
.C(n_13),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_465),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_470),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_13),
.B(n_487),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_472),
.C(n_483),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_492),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_493),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_486),
.C(n_491),
.Y(n_498)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_498),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_495),
.B(n_494),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_500),
.A2(n_499),
.B(n_13),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_501),
.Y(n_503)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_503),
.Y(n_504)
);


endmodule