module fake_netlist_6_4766_n_5344 (n_992, n_1, n_801, n_1234, n_1199, n_741, n_1027, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1038, n_578, n_1003, n_365, n_168, n_1237, n_1061, n_77, n_783, n_798, n_188, n_509, n_245, n_1209, n_677, n_805, n_1151, n_396, n_350, n_78, n_442, n_480, n_142, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_893, n_1099, n_1192, n_471, n_424, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_200, n_447, n_1172, n_852, n_71, n_229, n_1078, n_250, n_544, n_1140, n_35, n_836, n_375, n_522, n_1261, n_945, n_1143, n_1232, n_616, n_658, n_1119, n_428, n_641, n_822, n_693, n_1056, n_758, n_516, n_1163, n_1180, n_943, n_491, n_42, n_772, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_343, n_953, n_1094, n_494, n_539, n_493, n_155, n_45, n_454, n_638, n_1211, n_381, n_887, n_112, n_713, n_126, n_58, n_976, n_224, n_48, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_14, n_659, n_407, n_913, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_44, n_163, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_577, n_166, n_619, n_521, n_572, n_395, n_813, n_323, n_606, n_818, n_1123, n_92, n_513, n_645, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_219, n_264, n_263, n_1162, n_860, n_788, n_939, n_821, n_938, n_1068, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_117, n_175, n_322, n_993, n_689, n_354, n_134, n_547, n_558, n_1064, n_634, n_136, n_966, n_764, n_692, n_733, n_1233, n_487, n_241, n_30, n_1107, n_1014, n_882, n_586, n_423, n_318, n_1111, n_715, n_1251, n_88, n_530, n_277, n_618, n_199, n_1167, n_674, n_871, n_922, n_268, n_210, n_1069, n_5, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_429, n_1012, n_195, n_780, n_675, n_903, n_286, n_254, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_816, n_1157, n_1188, n_877, n_604, n_825, n_728, n_1063, n_26, n_55, n_267, n_1124, n_515, n_598, n_696, n_961, n_437, n_1082, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_949, n_678, n_283, n_91, n_507, n_968, n_909, n_881, n_1008, n_760, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_304, n_694, n_125, n_297, n_595, n_627, n_524, n_342, n_1044, n_449, n_131, n_1208, n_1164, n_1072, n_495, n_815, n_1100, n_585, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_615, n_1249, n_59, n_1127, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_826, n_872, n_1139, n_86, n_104, n_718, n_1018, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_413, n_791, n_510, n_837, n_79, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_581, n_765, n_432, n_987, n_631, n_720, n_153, n_842, n_156, n_145, n_843, n_656, n_989, n_797, n_1246, n_899, n_189, n_738, n_1035, n_294, n_499, n_705, n_11, n_1004, n_1176, n_1022, n_614, n_529, n_425, n_684, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_648, n_657, n_1049, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_777, n_272, n_526, n_1183, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_18, n_154, n_1178, n_98, n_1073, n_1000, n_796, n_252, n_1195, n_184, n_552, n_216, n_912, n_745, n_1142, n_716, n_623, n_1048, n_1201, n_884, n_731, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_66, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_589, n_819, n_767, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_399, n_124, n_211, n_231, n_40, n_505, n_319, n_537, n_311, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_386, n_1220, n_556, n_162, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1053, n_416, n_520, n_418, n_1093, n_113, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_217, n_518, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_90, n_54, n_488, n_497, n_773, n_920, n_99, n_13, n_1224, n_1135, n_1169, n_1179, n_401, n_324, n_335, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_36, n_983, n_427, n_496, n_906, n_688, n_1077, n_351, n_259, n_177, n_385, n_858, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1134, n_410, n_1129, n_554, n_602, n_664, n_171, n_169, n_435, n_793, n_326, n_587, n_580, n_762, n_1030, n_1202, n_465, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_485, n_67, n_443, n_892, n_768, n_421, n_238, n_1095, n_202, n_597, n_280, n_1187, n_610, n_1024, n_198, n_179, n_248, n_517, n_667, n_1206, n_621, n_1037, n_1115, n_750, n_901, n_468, n_923, n_504, n_183, n_1015, n_466, n_1057, n_603, n_991, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_39, n_73, n_785, n_746, n_609, n_101, n_167, n_127, n_1168, n_1216, n_133, n_96, n_302, n_380, n_137, n_20, n_1190, n_397, n_122, n_34, n_218, n_1213, n_70, n_172, n_239, n_97, n_782, n_490, n_220, n_809, n_1043, n_986, n_80, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_662, n_374, n_1152, n_450, n_921, n_711, n_579, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_258, n_456, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_936, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_420, n_394, n_164, n_23, n_942, n_543, n_1225, n_325, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_76, n_548, n_94, n_282, n_833, n_523, n_707, n_345, n_799, n_1155, n_139, n_41, n_273, n_787, n_1146, n_159, n_1086, n_1066, n_157, n_550, n_275, n_652, n_560, n_1241, n_569, n_737, n_1235, n_1229, n_306, n_21, n_346, n_3, n_1029, n_790, n_138, n_1210, n_49, n_299, n_1248, n_902, n_333, n_1047, n_431, n_24, n_459, n_502, n_672, n_1257, n_285, n_85, n_655, n_706, n_1045, n_786, n_1236, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_660, n_438, n_1200, n_479, n_869, n_1154, n_1113, n_646, n_528, n_391, n_1098, n_817, n_262, n_187, n_897, n_846, n_841, n_1001, n_508, n_1050, n_1177, n_332, n_1150, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_855, n_52, n_591, n_256, n_853, n_440, n_695, n_875, n_209, n_367, n_680, n_661, n_278, n_1256, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1217, n_751, n_749, n_310, n_969, n_988, n_1065, n_84, n_1255, n_568, n_143, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_739, n_400, n_955, n_337, n_214, n_246, n_1097, n_935, n_781, n_789, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_555, n_389, n_814, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1105, n_721, n_742, n_535, n_691, n_372, n_111, n_314, n_378, n_1196, n_377, n_863, n_601, n_338, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_119, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1205, n_1258, n_174, n_1173, n_525, n_1116, n_611, n_1219, n_8, n_1174, n_1016, n_795, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_930, n_888, n_1112, n_234, n_910, n_911, n_82, n_27, n_236, n_653, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_779, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_366, n_103, n_1109, n_185, n_712, n_348, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_470, n_475, n_924, n_298, n_492, n_1149, n_265, n_1184, n_228, n_719, n_455, n_363, n_1090, n_592, n_829, n_1156, n_393, n_984, n_503, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_981, n_714, n_291, n_1144, n_357, n_985, n_481, n_997, n_802, n_561, n_33, n_980, n_1198, n_436, n_116, n_409, n_1244, n_240, n_756, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_583, n_249, n_201, n_1039, n_1034, n_1158, n_754, n_941, n_975, n_1031, n_115, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1055, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_588, n_225, n_1260, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1006, n_373, n_87, n_257, n_730, n_670, n_203, n_207, n_1089, n_205, n_1242, n_681, n_1226, n_412, n_640, n_81, n_965, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_457, n_364, n_629, n_900, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_1259, n_192, n_51, n_649, n_1240, n_5344);

input n_992;
input n_1;
input n_801;
input n_1234;
input n_1199;
input n_741;
input n_1027;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1038;
input n_578;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_77;
input n_783;
input n_798;
input n_188;
input n_509;
input n_245;
input n_1209;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_442;
input n_480;
input n_142;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_893;
input n_1099;
input n_1192;
input n_471;
input n_424;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_35;
input n_836;
input n_375;
input n_522;
input n_1261;
input n_945;
input n_1143;
input n_1232;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_758;
input n_516;
input n_1163;
input n_1180;
input n_943;
input n_491;
input n_42;
input n_772;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_343;
input n_953;
input n_1094;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_638;
input n_1211;
input n_381;
input n_887;
input n_112;
input n_713;
input n_126;
input n_58;
input n_976;
input n_224;
input n_48;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_14;
input n_659;
input n_407;
input n_913;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_44;
input n_163;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_577;
input n_166;
input n_619;
input n_521;
input n_572;
input n_395;
input n_813;
input n_323;
input n_606;
input n_818;
input n_1123;
input n_92;
input n_513;
input n_645;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_788;
input n_939;
input n_821;
input n_938;
input n_1068;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_134;
input n_547;
input n_558;
input n_1064;
input n_634;
input n_136;
input n_966;
input n_764;
input n_692;
input n_733;
input n_1233;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_882;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_88;
input n_530;
input n_277;
input n_618;
input n_199;
input n_1167;
input n_674;
input n_871;
input n_922;
input n_268;
input n_210;
input n_1069;
input n_5;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_286;
input n_254;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_816;
input n_1157;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_515;
input n_598;
input n_696;
input n_961;
input n_437;
input n_1082;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_949;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_881;
input n_1008;
input n_760;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_304;
input n_694;
input n_125;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_1044;
input n_449;
input n_131;
input n_1208;
input n_1164;
input n_1072;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_615;
input n_1249;
input n_59;
input n_1127;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_826;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_581;
input n_765;
input n_432;
input n_987;
input n_631;
input n_720;
input n_153;
input n_842;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_797;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1035;
input n_294;
input n_499;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_648;
input n_657;
input n_1049;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_777;
input n_272;
input n_526;
input n_1183;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_18;
input n_154;
input n_1178;
input n_98;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_184;
input n_552;
input n_216;
input n_912;
input n_745;
input n_1142;
input n_716;
input n_623;
input n_1048;
input n_1201;
input n_884;
input n_731;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_66;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_589;
input n_819;
input n_767;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_399;
input n_124;
input n_211;
input n_231;
input n_40;
input n_505;
input n_319;
input n_537;
input n_311;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_217;
input n_518;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_90;
input n_54;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_13;
input n_1224;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_335;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_36;
input n_983;
input n_427;
input n_496;
input n_906;
input n_688;
input n_1077;
input n_351;
input n_259;
input n_177;
input n_385;
input n_858;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_664;
input n_171;
input n_169;
input n_435;
input n_793;
input n_326;
input n_587;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_485;
input n_67;
input n_443;
input n_892;
input n_768;
input n_421;
input n_238;
input n_1095;
input n_202;
input n_597;
input n_280;
input n_1187;
input n_610;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1115;
input n_750;
input n_901;
input n_468;
input n_923;
input n_504;
input n_183;
input n_1015;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_39;
input n_73;
input n_785;
input n_746;
input n_609;
input n_101;
input n_167;
input n_127;
input n_1168;
input n_1216;
input n_133;
input n_96;
input n_302;
input n_380;
input n_137;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_218;
input n_1213;
input n_70;
input n_172;
input n_239;
input n_97;
input n_782;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_986;
input n_80;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_711;
input n_579;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_258;
input n_456;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_936;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_420;
input n_394;
input n_164;
input n_23;
input n_942;
input n_543;
input n_1225;
input n_325;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_76;
input n_548;
input n_94;
input n_282;
input n_833;
input n_523;
input n_707;
input n_345;
input n_799;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_787;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1241;
input n_569;
input n_737;
input n_1235;
input n_1229;
input n_306;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_790;
input n_138;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_333;
input n_1047;
input n_431;
input n_24;
input n_459;
input n_502;
input n_672;
input n_1257;
input n_285;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_786;
input n_1236;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_660;
input n_438;
input n_1200;
input n_479;
input n_869;
input n_1154;
input n_1113;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1001;
input n_508;
input n_1050;
input n_1177;
input n_332;
input n_1150;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_855;
input n_52;
input n_591;
input n_256;
input n_853;
input n_440;
input n_695;
input n_875;
input n_209;
input n_367;
input n_680;
input n_661;
input n_278;
input n_1256;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_1255;
input n_568;
input n_143;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_739;
input n_400;
input n_955;
input n_337;
input n_214;
input n_246;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_555;
input n_389;
input n_814;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1105;
input n_721;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_378;
input n_1196;
input n_377;
input n_863;
input n_601;
input n_338;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_119;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1205;
input n_1258;
input n_174;
input n_1173;
input n_525;
input n_1116;
input n_611;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_795;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_911;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_779;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_366;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_455;
input n_363;
input n_1090;
input n_592;
input n_829;
input n_1156;
input n_393;
input n_984;
input n_503;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_981;
input n_714;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1198;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_240;
input n_756;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1034;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1055;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1006;
input n_373;
input n_87;
input n_257;
input n_730;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_412;
input n_640;
input n_81;
input n_965;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_457;
input n_364;
input n_629;
input n_900;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_1259;
input n_192;
input n_51;
input n_649;
input n_1240;

output n_5344;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_1351;
wire n_5254;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_3089;
wire n_4978;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5332;
wire n_2004;
wire n_4814;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_2764;
wire n_2895;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_5183;
wire n_2145;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1512;
wire n_1451;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_3179;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_4345;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_4528;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_5035;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_1955;
wire n_1791;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_4189;
wire n_3817;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_4512;
wire n_1378;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_5124;
wire n_3951;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_3027;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2020;
wire n_1643;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1461;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_4027;
wire n_3154;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1570;
wire n_1702;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1574;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_5335;
wire n_3444;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_3017;
wire n_1890;
wire n_2477;
wire n_1805;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_3266;
wire n_3574;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_4504;
wire n_3844;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_5248;
wire n_1708;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1511;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_4047;
wire n_3413;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_3725;
wire n_3933;
wire n_2311;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_2271;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_3431;
wire n_1767;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_2954;
wire n_2728;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_3442;
wire n_1880;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_5087;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_1959;
wire n_5257;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_2338;
wire n_3324;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_5282;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1951;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_4404;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_2315;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_3250;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1683;
wire n_1916;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_4016;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2808;
wire n_2037;
wire n_4567;
wire n_5150;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_2390;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_4143;
wire n_4170;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_3515;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_4910;
wire n_3083;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_4521;
wire n_1566;
wire n_3204;
wire n_4920;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_4730;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2256;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_2806;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_3568;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1530;
wire n_4745;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_3599;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_4800;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_3326;
wire n_2036;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_3805;
wire n_1990;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_4097;
wire n_1666;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_3636;
wire n_2327;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_2755;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1692;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_2699;
wire n_1828;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_1405;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_2141;
wire n_5316;
wire n_3930;
wire n_4943;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_2021;
wire n_4942;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_3157;
wire n_4841;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_5320;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_2045;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_2566;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_2042;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_4089;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_4865;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1819;
wire n_3555;
wire n_3155;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_2336;
wire n_2521;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_3822;
wire n_4163;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_4372;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_4673;
wire n_2519;
wire n_3415;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_4019;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_3144;
wire n_3244;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2357;
wire n_2025;
wire n_4654;
wire n_3640;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_2278;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_2704;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_1794;
wire n_4493;
wire n_4924;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_2066;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1327;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_2380;
wire n_4786;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_3493;
wire n_3774;
wire n_2910;
wire n_3268;
wire n_1785;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_2287;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_3334;
wire n_5097;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_2600;
wire n_3508;
wire n_4353;
wire n_4787;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_2440;
wire n_3521;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_2909;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1185),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_357),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_221),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1075),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_777),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_789),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_172),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1222),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_457),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_236),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_773),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_786),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_407),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1140),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_432),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1153),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1229),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1240),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_391),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_607),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_195),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_367),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1019),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_835),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1008),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_507),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1195),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_734),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1035),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_471),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_961),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_980),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_903),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_991),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1116),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_295),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_130),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1091),
.Y(n_1299)
);

CKINVDCx14_ASAP7_75t_R g1300 ( 
.A(n_149),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1122),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_776),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_343),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_775),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_962),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1214),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_929),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1000),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1182),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_15),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_238),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1137),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_270),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1226),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_983),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_689),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_14),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1179),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_722),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_998),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1087),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1032),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_107),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_691),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_121),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1154),
.Y(n_1326)
);

CKINVDCx14_ASAP7_75t_R g1327 ( 
.A(n_879),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1251),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_764),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_914),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_566),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_185),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1065),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_111),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_986),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_242),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_249),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_132),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_8),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_936),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_637),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_726),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_42),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_819),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_999),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1183),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_596),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_884),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_292),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_42),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1096),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1152),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_839),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_241),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_813),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_920),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1080),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1181),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1077),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_110),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_59),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1191),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_808),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_997),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_372),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1024),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_972),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1125),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1236),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_555),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1042),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_365),
.Y(n_1372)
);

CKINVDCx14_ASAP7_75t_R g1373 ( 
.A(n_663),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_459),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1151),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_536),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_706),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_549),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_288),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1201),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1107),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1033),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_960),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_381),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1130),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_786),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1259),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_79),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_840),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_842),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_959),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_941),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_951),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_928),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1009),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1110),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_733),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1081),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_261),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1218),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_839),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_360),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1090),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_26),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1217),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1118),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1166),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_880),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1172),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1002),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_503),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_979),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_441),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1034),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_27),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1020),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_191),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_946),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_963),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_121),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_132),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_782),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_210),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_750),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_932),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_804),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_511),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1221),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_937),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1207),
.Y(n_1430)
);

BUFx10_ASAP7_75t_L g1431 ( 
.A(n_1228),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_698),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_598),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_183),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1244),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_719),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_513),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_184),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_62),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1027),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_214),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_989),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_508),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_636),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_24),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_32),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_417),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_911),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_62),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1039),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_958),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_968),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1061),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_270),
.Y(n_1454)
);

BUFx10_ASAP7_75t_L g1455 ( 
.A(n_174),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1089),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_641),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_409),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_37),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_645),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_941),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1243),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_73),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_783),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1015),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_443),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_117),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1176),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_863),
.Y(n_1469)
);

BUFx10_ASAP7_75t_L g1470 ( 
.A(n_1170),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_838),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_234),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1076),
.Y(n_1473)
);

CKINVDCx16_ASAP7_75t_R g1474 ( 
.A(n_1131),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_981),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_87),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_214),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_721),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_321),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_807),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_943),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_944),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_229),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_17),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1088),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_857),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_449),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1252),
.Y(n_1488)
);

BUFx5_ASAP7_75t_L g1489 ( 
.A(n_1101),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1213),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_600),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_855),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1053),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_952),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1121),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1049),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_254),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_397),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_587),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_343),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_752),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1031),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_166),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_126),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1112),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_91),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_123),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_514),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1094),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1138),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_554),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1012),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1205),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1111),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_233),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_193),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_597),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_174),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1219),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_576),
.Y(n_1520)
);

BUFx10_ASAP7_75t_L g1521 ( 
.A(n_542),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_238),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1123),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_526),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1008),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1197),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_303),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1126),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1160),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_1158),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1250),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1150),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1254),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1168),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_632),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_905),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_542),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_465),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1104),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_378),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_761),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1178),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1142),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_649),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1189),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_683),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_970),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_638),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_30),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_862),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_56),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_597),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1040),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_686),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_237),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_990),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1256),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_832),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_807),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1010),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_466),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_334),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_623),
.Y(n_1563)
);

BUFx2_ASAP7_75t_SL g1564 ( 
.A(n_923),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_927),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_996),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_141),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1139),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1011),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_82),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1188),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_879),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_167),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_614),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_362),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_574),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_973),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_810),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_754),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_933),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_955),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_160),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_548),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_16),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_94),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1233),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1102),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_658),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_926),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_39),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_995),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_545),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1200),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_634),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_830),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1212),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_974),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1099),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_853),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_795),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1128),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_759),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1194),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_671),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_736),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_477),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_141),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_961),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1144),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_655),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1261),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_364),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_504),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_978),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_278),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_598),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_861),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_686),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1136),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_257),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1103),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_664),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_256),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_922),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_142),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_985),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_991),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1167),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1159),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_432),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_399),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1155),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_541),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1235),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_339),
.Y(n_1635)
);

INVxp33_ASAP7_75t_R g1636 ( 
.A(n_49),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1120),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_958),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1257),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_950),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_382),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_587),
.Y(n_1642)
);

CKINVDCx14_ASAP7_75t_R g1643 ( 
.A(n_199),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_340),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_396),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_600),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_20),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_409),
.Y(n_1648)
);

BUFx10_ASAP7_75t_L g1649 ( 
.A(n_473),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_678),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_927),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_250),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_954),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_428),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_219),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_643),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_315),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_329),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_849),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1239),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_341),
.Y(n_1661)
);

CKINVDCx14_ASAP7_75t_R g1662 ( 
.A(n_813),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_229),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_755),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_5),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_956),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_801),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1097),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1210),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1174),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_701),
.Y(n_1671)
);

BUFx10_ASAP7_75t_L g1672 ( 
.A(n_387),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_282),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_675),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1068),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_695),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_162),
.Y(n_1677)
);

BUFx10_ASAP7_75t_L g1678 ( 
.A(n_1211),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1260),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1227),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1215),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_422),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_769),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_463),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1001),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_582),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_976),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1117),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1098),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_592),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_658),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_566),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1082),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1109),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_212),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_539),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_812),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_948),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_849),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_628),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_501),
.Y(n_1701)
);

BUFx5_ASAP7_75t_L g1702 ( 
.A(n_1225),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_45),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1148),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_498),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_265),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_66),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_953),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1193),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1079),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_414),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_855),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1202),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1145),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_468),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1149),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_659),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1164),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_462),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1134),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_474),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_793),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1007),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1074),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1085),
.Y(n_1725)
);

BUFx5_ASAP7_75t_L g1726 ( 
.A(n_881),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_965),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1133),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_498),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_279),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_648),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_113),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_925),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_971),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_461),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_960),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_946),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_147),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1196),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_911),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_607),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_184),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_81),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_593),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_144),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_188),
.Y(n_1746)
);

BUFx10_ASAP7_75t_L g1747 ( 
.A(n_12),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_676),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1105),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_957),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_661),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_375),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1187),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_183),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_279),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_437),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_969),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_893),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_967),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_900),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_676),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1237),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1253),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_427),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1161),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_640),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_378),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1177),
.Y(n_1768)
);

BUFx8_ASAP7_75t_SL g1769 ( 
.A(n_501),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_240),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1156),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_556),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_903),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_935),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_988),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_371),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_389),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_160),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1006),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_873),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1245),
.Y(n_1781)
);

BUFx10_ASAP7_75t_L g1782 ( 
.A(n_965),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_694),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1247),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1029),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_290),
.Y(n_1786)
);

BUFx10_ASAP7_75t_L g1787 ( 
.A(n_868),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_408),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_1132),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1046),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_668),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_708),
.Y(n_1792)
);

BUFx10_ASAP7_75t_L g1793 ( 
.A(n_838),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_843),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1190),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_572),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1175),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_804),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_655),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1163),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1186),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1003),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_688),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_399),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_363),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_208),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1206),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_404),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_803),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_939),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1004),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_949),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1083),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1249),
.Y(n_1814)
);

INVx2_ASAP7_75t_SL g1815 ( 
.A(n_947),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_6),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1124),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1129),
.Y(n_1818)
);

CKINVDCx16_ASAP7_75t_R g1819 ( 
.A(n_915),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_603),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_489),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_522),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_478),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_691),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_400),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_549),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_420),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_355),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_202),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1157),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_406),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_81),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_162),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_993),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_771),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_530),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_291),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_792),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_564),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_978),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_715),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_321),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_125),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_294),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_390),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_888),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1043),
.Y(n_1847)
);

BUFx10_ASAP7_75t_L g1848 ( 
.A(n_1162),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1146),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_826),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_657),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_982),
.Y(n_1852)
);

BUFx10_ASAP7_75t_L g1853 ( 
.A(n_227),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_923),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1192),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_609),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1047),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1199),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_47),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_940),
.Y(n_1860)
);

CKINVDCx16_ASAP7_75t_R g1861 ( 
.A(n_865),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_318),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1135),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_822),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1242),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_136),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_147),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_894),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1095),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_0),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_443),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1203),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_654),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1086),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_313),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1198),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_977),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_16),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_395),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_975),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_71),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_649),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_288),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_671),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_78),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_735),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_916),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_893),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1078),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_318),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_479),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_936),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1108),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_528),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_714),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_614),
.B(n_966),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_712),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_948),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_924),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_113),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1171),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1017),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_302),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_468),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_303),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1070),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_458),
.Y(n_1907)
);

BUFx10_ASAP7_75t_L g1908 ( 
.A(n_1026),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_299),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_334),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1223),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_492),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1069),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1234),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_430),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_513),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_525),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1141),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_826),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1180),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1184),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_921),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1204),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_701),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_987),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_931),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_416),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1084),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_367),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_299),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1127),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_7),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1062),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1030),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_934),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1005),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_172),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_351),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_317),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_129),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1216),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1147),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_26),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_994),
.Y(n_1944)
);

CKINVDCx20_ASAP7_75t_R g1945 ( 
.A(n_1113),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_28),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_726),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_212),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_144),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_494),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_591),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_471),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_429),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1114),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_942),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_127),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_216),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_352),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_336),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_992),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1092),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_929),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_463),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_493),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_485),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1208),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_306),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_641),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_872),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_553),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_531),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_827),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_930),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_964),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_837),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_156),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_798),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_441),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_624),
.Y(n_1979)
);

CKINVDCx14_ASAP7_75t_R g1980 ( 
.A(n_918),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_99),
.Y(n_1981)
);

INVxp67_ASAP7_75t_SL g1982 ( 
.A(n_371),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_905),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_792),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1169),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1143),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1173),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_234),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_574),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_400),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_672),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_866),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_670),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_938),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_642),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_945),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_984),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1064),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_100),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1209),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_272),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1100),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_227),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_123),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_683),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_733),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1115),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_326),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1230),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_527),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_986),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_397),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_687),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_875),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_781),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1009),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1241),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_416),
.Y(n_2018)
);

CKINVDCx20_ASAP7_75t_R g2019 ( 
.A(n_546),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1231),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_624),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1119),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_5),
.Y(n_2023)
);

CKINVDCx20_ASAP7_75t_R g2024 ( 
.A(n_631),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1106),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_287),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_705),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_429),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1093),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_647),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1071),
.Y(n_2031)
);

BUFx5_ASAP7_75t_L g2032 ( 
.A(n_651),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1165),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_173),
.Y(n_2034)
);

BUFx10_ASAP7_75t_L g2035 ( 
.A(n_939),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_573),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1246),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1238),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_871),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1248),
.Y(n_2040)
);

BUFx10_ASAP7_75t_L g2041 ( 
.A(n_523),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_236),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_837),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_631),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1232),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1050),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_483),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_40),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_52),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_20),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1258),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_260),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_476),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1255),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_206),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_659),
.Y(n_2056)
);

CKINVDCx20_ASAP7_75t_R g2057 ( 
.A(n_401),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_880),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_667),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_484),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_796),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_1220),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_693),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1224),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1726),
.Y(n_2065)
);

INVxp33_ASAP7_75t_L g2066 ( 
.A(n_1311),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1769),
.Y(n_2067)
);

BUFx2_ASAP7_75t_SL g2068 ( 
.A(n_1381),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1431),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_1542),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1726),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1348),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1726),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1435),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1726),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1726),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2032),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2032),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2032),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1269),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1402),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2032),
.Y(n_2082)
);

INVxp33_ASAP7_75t_L g2083 ( 
.A(n_1379),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2032),
.Y(n_2084)
);

INVx2_ASAP7_75t_SL g2085 ( 
.A(n_1391),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1275),
.Y(n_2086)
);

INVxp33_ASAP7_75t_L g2087 ( 
.A(n_1420),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1402),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1402),
.Y(n_2089)
);

INVxp33_ASAP7_75t_L g2090 ( 
.A(n_1479),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1487),
.Y(n_2091)
);

INVxp33_ASAP7_75t_SL g2092 ( 
.A(n_1585),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1487),
.Y(n_2093)
);

CKINVDCx16_ASAP7_75t_R g2094 ( 
.A(n_1340),
.Y(n_2094)
);

CKINVDCx16_ASAP7_75t_R g2095 ( 
.A(n_1451),
.Y(n_2095)
);

CKINVDCx20_ASAP7_75t_R g2096 ( 
.A(n_1611),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1277),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_1484),
.Y(n_2098)
);

INVxp33_ASAP7_75t_SL g2099 ( 
.A(n_1667),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_1565),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1487),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1278),
.Y(n_2102)
);

INVxp67_ASAP7_75t_SL g2103 ( 
.A(n_1262),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1582),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1582),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1582),
.Y(n_2106)
);

INVxp33_ASAP7_75t_SL g2107 ( 
.A(n_2056),
.Y(n_2107)
);

CKINVDCx16_ASAP7_75t_R g2108 ( 
.A(n_1497),
.Y(n_2108)
);

CKINVDCx16_ASAP7_75t_R g2109 ( 
.A(n_1551),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1602),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1602),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1296),
.Y(n_2112)
);

INVxp33_ASAP7_75t_L g2113 ( 
.A(n_1578),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1602),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_1593),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1706),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1706),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1706),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1711),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1299),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1711),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1711),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_1306),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1712),
.Y(n_2124)
);

BUFx3_ASAP7_75t_L g2125 ( 
.A(n_1431),
.Y(n_2125)
);

CKINVDCx16_ASAP7_75t_R g2126 ( 
.A(n_1819),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1712),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1712),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_1284),
.B(n_1),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1783),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1783),
.Y(n_2131)
);

NOR2xp67_ASAP7_75t_L g2132 ( 
.A(n_1896),
.B(n_0),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1783),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_1650),
.Y(n_2134)
);

INVxp33_ASAP7_75t_SL g2135 ( 
.A(n_1671),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1835),
.Y(n_2136)
);

CKINVDCx20_ASAP7_75t_R g2137 ( 
.A(n_1668),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1835),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1835),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1884),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_1834),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1309),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1318),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1884),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1845),
.Y(n_2145)
);

INVxp33_ASAP7_75t_SL g2146 ( 
.A(n_1864),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1884),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1994),
.Y(n_2148)
);

INVxp33_ASAP7_75t_SL g2149 ( 
.A(n_1975),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1321),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1326),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1994),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_1994),
.Y(n_2153)
);

INVxp67_ASAP7_75t_SL g2154 ( 
.A(n_2020),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1328),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1489),
.Y(n_2156)
);

BUFx10_ASAP7_75t_L g2157 ( 
.A(n_1266),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1283),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1441),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1478),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1516),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1541),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1391),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1659),
.Y(n_2164)
);

INVxp33_ASAP7_75t_L g2165 ( 
.A(n_2028),
.Y(n_2165)
);

CKINVDCx16_ASAP7_75t_R g2166 ( 
.A(n_1861),
.Y(n_2166)
);

INVxp67_ASAP7_75t_SL g2167 ( 
.A(n_1533),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1661),
.Y(n_2168)
);

CKINVDCx20_ASAP7_75t_R g2169 ( 
.A(n_1789),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1333),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1352),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1489),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1673),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1357),
.Y(n_2174)
);

CKINVDCx20_ASAP7_75t_R g2175 ( 
.A(n_1801),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1686),
.Y(n_2176)
);

NOR2xp67_ASAP7_75t_L g2177 ( 
.A(n_1386),
.B(n_1),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1359),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1489),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1362),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1489),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1489),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2063),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1263),
.Y(n_2184)
);

INVxp33_ASAP7_75t_SL g2185 ( 
.A(n_1267),
.Y(n_2185)
);

INVxp67_ASAP7_75t_SL g2186 ( 
.A(n_1279),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2052),
.Y(n_2187)
);

CKINVDCx20_ASAP7_75t_R g2188 ( 
.A(n_1865),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1271),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1272),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1273),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1281),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1291),
.Y(n_2193)
);

INVxp33_ASAP7_75t_SL g2194 ( 
.A(n_1268),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1305),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1310),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1315),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1324),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1330),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1334),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1347),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1349),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1353),
.Y(n_2203)
);

INVxp67_ASAP7_75t_SL g2204 ( 
.A(n_1290),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_1300),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1354),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1361),
.Y(n_2207)
);

CKINVDCx16_ASAP7_75t_R g2208 ( 
.A(n_1474),
.Y(n_2208)
);

INVxp33_ASAP7_75t_L g2209 ( 
.A(n_1365),
.Y(n_2209)
);

INVxp67_ASAP7_75t_SL g2210 ( 
.A(n_1495),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1367),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1372),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1376),
.Y(n_2213)
);

INVxp67_ASAP7_75t_SL g2214 ( 
.A(n_1637),
.Y(n_2214)
);

INVxp67_ASAP7_75t_SL g2215 ( 
.A(n_1728),
.Y(n_2215)
);

INVxp33_ASAP7_75t_SL g2216 ( 
.A(n_1276),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1702),
.Y(n_2217)
);

CKINVDCx20_ASAP7_75t_R g2218 ( 
.A(n_1942),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1384),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1393),
.Y(n_2220)
);

CKINVDCx16_ASAP7_75t_R g2221 ( 
.A(n_1327),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1395),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1397),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1264),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1415),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1426),
.Y(n_2226)
);

INVxp67_ASAP7_75t_SL g2227 ( 
.A(n_1918),
.Y(n_2227)
);

INVxp67_ASAP7_75t_SL g2228 ( 
.A(n_1288),
.Y(n_2228)
);

OA21x2_ASAP7_75t_L g2229 ( 
.A1(n_2065),
.A2(n_1314),
.B(n_1301),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2089),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2205),
.B(n_1373),
.Y(n_2231)
);

BUFx3_ASAP7_75t_L g2232 ( 
.A(n_2158),
.Y(n_2232)
);

OAI21x1_ASAP7_75t_L g2233 ( 
.A1(n_2156),
.A2(n_1312),
.B(n_1265),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_2069),
.B(n_1704),
.Y(n_2234)
);

INVx5_ASAP7_75t_L g2235 ( 
.A(n_2157),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_2081),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2091),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2127),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2186),
.B(n_1643),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2094),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2144),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2185),
.B(n_1662),
.Y(n_2242)
);

INVx5_ASAP7_75t_L g2243 ( 
.A(n_2157),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2147),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2125),
.B(n_1724),
.Y(n_2245)
);

AOI22x1_ASAP7_75t_SL g2246 ( 
.A1(n_2070),
.A2(n_1285),
.B1(n_1289),
.B2(n_1270),
.Y(n_2246)
);

OAI22x1_ASAP7_75t_R g2247 ( 
.A1(n_2096),
.A2(n_1298),
.B1(n_1303),
.B2(n_1297),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2088),
.Y(n_2248)
);

INVx2_ASAP7_75t_SL g2249 ( 
.A(n_2085),
.Y(n_2249)
);

BUFx8_ASAP7_75t_L g2250 ( 
.A(n_2145),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2194),
.B(n_1980),
.Y(n_2251)
);

BUFx8_ASAP7_75t_L g2252 ( 
.A(n_2163),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2074),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2074),
.Y(n_2254)
);

BUFx12f_ASAP7_75t_L g2255 ( 
.A(n_2067),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_2074),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2204),
.B(n_1470),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2081),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2153),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2153),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2080),
.B(n_1450),
.Y(n_2261)
);

OAI21x1_ASAP7_75t_L g2262 ( 
.A1(n_2172),
.A2(n_1430),
.B(n_1406),
.Y(n_2262)
);

AOI22x1_ASAP7_75t_SL g2263 ( 
.A1(n_2137),
.A2(n_1364),
.B1(n_1383),
.B2(n_1307),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2135),
.A2(n_1945),
.B1(n_1982),
.B2(n_1280),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2093),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2210),
.B(n_1470),
.Y(n_2266)
);

INVx4_ASAP7_75t_L g2267 ( 
.A(n_2086),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2097),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2101),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2104),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2102),
.B(n_1490),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2105),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2167),
.B(n_1813),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2106),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2095),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2110),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2214),
.B(n_1768),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_2159),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2108),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2111),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2146),
.A2(n_1287),
.B1(n_1292),
.B2(n_1286),
.Y(n_2281)
);

INVx5_ASAP7_75t_L g2282 ( 
.A(n_2221),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2112),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_2160),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2120),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2114),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2116),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_2224),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2117),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2118),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2123),
.B(n_2062),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2119),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2142),
.B(n_1465),
.Y(n_2293)
);

BUFx8_ASAP7_75t_L g2294 ( 
.A(n_2161),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2121),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2149),
.A2(n_1302),
.B1(n_1304),
.B2(n_1293),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2092),
.A2(n_1657),
.B1(n_1936),
.B2(n_1584),
.Y(n_2297)
);

AOI22x1_ASAP7_75t_SL g2298 ( 
.A1(n_2169),
.A2(n_1491),
.B1(n_1506),
.B2(n_1472),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2143),
.B(n_1488),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2122),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_2124),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2128),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2130),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2150),
.B(n_1502),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2131),
.Y(n_2305)
);

INVx3_ASAP7_75t_L g2306 ( 
.A(n_2224),
.Y(n_2306)
);

OAI21x1_ASAP7_75t_L g2307 ( 
.A1(n_2179),
.A2(n_1601),
.B(n_1543),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2133),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2136),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2138),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2139),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2099),
.A2(n_1313),
.B1(n_1319),
.B2(n_1317),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2140),
.Y(n_2313)
);

INVx3_ASAP7_75t_L g2314 ( 
.A(n_2148),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2152),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_2151),
.Y(n_2316)
);

OAI21x1_ASAP7_75t_L g2317 ( 
.A1(n_2181),
.A2(n_2217),
.B(n_2182),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2071),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2215),
.B(n_1322),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_2183),
.Y(n_2320)
);

INVx5_ASAP7_75t_L g2321 ( 
.A(n_2109),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2107),
.A2(n_1320),
.B1(n_1325),
.B2(n_1323),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_L g2323 ( 
.A(n_2073),
.B(n_1346),
.Y(n_2323)
);

INVx4_ASAP7_75t_L g2324 ( 
.A(n_2155),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2075),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_2170),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_2184),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2076),
.Y(n_2328)
);

CKINVDCx6p67_ASAP7_75t_R g2329 ( 
.A(n_2126),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_2187),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_2171),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2162),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2227),
.B(n_2103),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2216),
.B(n_2174),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2178),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2077),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_2180),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2078),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2115),
.B(n_1530),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2189),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2208),
.B(n_1530),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2079),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2082),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_2190),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2166),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2084),
.Y(n_2346)
);

INVx5_ASAP7_75t_L g2347 ( 
.A(n_2113),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2191),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2134),
.A2(n_1331),
.B1(n_1335),
.B2(n_1332),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2154),
.B(n_2072),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2192),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2193),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2195),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2228),
.B(n_1771),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2164),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2098),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2165),
.B(n_1678),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2066),
.B(n_1678),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2168),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2100),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2196),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2129),
.B(n_1351),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2197),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2141),
.B(n_1295),
.Y(n_2364)
);

BUFx8_ASAP7_75t_L g2365 ( 
.A(n_2173),
.Y(n_2365)
);

BUFx12f_ASAP7_75t_L g2366 ( 
.A(n_2068),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2198),
.Y(n_2367)
);

INVx5_ASAP7_75t_L g2368 ( 
.A(n_2083),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2199),
.Y(n_2369)
);

OA21x2_ASAP7_75t_L g2370 ( 
.A1(n_2200),
.A2(n_1382),
.B(n_1358),
.Y(n_2370)
);

BUFx3_ASAP7_75t_L g2371 ( 
.A(n_2176),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2201),
.Y(n_2372)
);

CKINVDCx8_ASAP7_75t_R g2373 ( 
.A(n_2175),
.Y(n_2373)
);

INVx2_ASAP7_75t_SL g2374 ( 
.A(n_2202),
.Y(n_2374)
);

BUFx8_ASAP7_75t_SL g2375 ( 
.A(n_2188),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2203),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2206),
.Y(n_2377)
);

INVx5_ASAP7_75t_L g2378 ( 
.A(n_2087),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2207),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2211),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2212),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2213),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2219),
.B(n_1863),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_2218),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2220),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2222),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2223),
.Y(n_2387)
);

BUFx2_ASAP7_75t_L g2388 ( 
.A(n_2225),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2090),
.B(n_1848),
.Y(n_2389)
);

OA21x2_ASAP7_75t_L g2390 ( 
.A1(n_2226),
.A2(n_1387),
.B(n_1385),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2177),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2209),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2132),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_2158),
.Y(n_2394)
);

OAI21x1_ASAP7_75t_L g2395 ( 
.A1(n_2156),
.A2(n_1941),
.B(n_1876),
.Y(n_2395)
);

AND2x6_ASAP7_75t_L g2396 ( 
.A(n_2129),
.B(n_1410),
.Y(n_2396)
);

BUFx8_ASAP7_75t_SL g2397 ( 
.A(n_2067),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_2080),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2089),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_2094),
.Y(n_2400)
);

INVx6_ASAP7_75t_L g2401 ( 
.A(n_2157),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2081),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2205),
.B(n_1396),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2205),
.B(n_1398),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2205),
.B(n_1409),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2089),
.Y(n_2406)
);

OAI21x1_ASAP7_75t_L g2407 ( 
.A1(n_2156),
.A2(n_2007),
.B(n_1453),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_2089),
.Y(n_2408)
);

INVx4_ASAP7_75t_L g2409 ( 
.A(n_2080),
.Y(n_2409)
);

INVx5_ASAP7_75t_L g2410 ( 
.A(n_2074),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2089),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2089),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_2080),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2081),
.Y(n_2414)
);

AND2x4_ASAP7_75t_L g2415 ( 
.A(n_2205),
.B(n_1440),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2080),
.B(n_1509),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_2069),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2080),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2089),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2089),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2089),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2069),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2205),
.B(n_1526),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2089),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2089),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_2080),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2205),
.B(n_1528),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2205),
.B(n_1848),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2081),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2205),
.B(n_1908),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2080),
.B(n_1531),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2080),
.B(n_1534),
.Y(n_2432)
);

INVx5_ASAP7_75t_L g2433 ( 
.A(n_2157),
.Y(n_2433)
);

HB1xp67_ASAP7_75t_L g2434 ( 
.A(n_2094),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2089),
.Y(n_2435)
);

INVx5_ASAP7_75t_L g2436 ( 
.A(n_2074),
.Y(n_2436)
);

INVx3_ASAP7_75t_L g2437 ( 
.A(n_2081),
.Y(n_2437)
);

AND2x6_ASAP7_75t_L g2438 ( 
.A(n_2129),
.B(n_1620),
.Y(n_2438)
);

INVx5_ASAP7_75t_L g2439 ( 
.A(n_2074),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_2080),
.Y(n_2440)
);

BUFx8_ASAP7_75t_L g2441 ( 
.A(n_2205),
.Y(n_2441)
);

INVx5_ASAP7_75t_L g2442 ( 
.A(n_2157),
.Y(n_2442)
);

OAI22x1_ASAP7_75t_SL g2443 ( 
.A1(n_2135),
.A2(n_1540),
.B1(n_1610),
.B2(n_1508),
.Y(n_2443)
);

BUFx12f_ASAP7_75t_L g2444 ( 
.A(n_2067),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2089),
.Y(n_2445)
);

OA21x2_ASAP7_75t_L g2446 ( 
.A1(n_2065),
.A2(n_1603),
.B(n_1598),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2089),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_2089),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2089),
.Y(n_2449)
);

AND2x4_ASAP7_75t_L g2450 ( 
.A(n_2205),
.B(n_1619),
.Y(n_2450)
);

OA21x2_ASAP7_75t_L g2451 ( 
.A1(n_2065),
.A2(n_1639),
.B(n_1628),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2089),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2089),
.Y(n_2453)
);

XNOR2xp5_ASAP7_75t_L g2454 ( 
.A(n_2070),
.B(n_1646),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2135),
.A2(n_1337),
.B1(n_1338),
.B2(n_1336),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2089),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2089),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2089),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2205),
.B(n_1669),
.Y(n_2459)
);

BUFx12f_ASAP7_75t_L g2460 ( 
.A(n_2067),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2080),
.B(n_1689),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2089),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2069),
.Y(n_2463)
);

OA21x2_ASAP7_75t_L g2464 ( 
.A1(n_2065),
.A2(n_1713),
.B(n_1709),
.Y(n_2464)
);

INVx3_ASAP7_75t_L g2465 ( 
.A(n_2081),
.Y(n_2465)
);

NOR2x1_ASAP7_75t_L g2466 ( 
.A(n_2069),
.B(n_1716),
.Y(n_2466)
);

BUFx12f_ASAP7_75t_L g2467 ( 
.A(n_2067),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2080),
.B(n_1718),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2089),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2205),
.B(n_1720),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2089),
.Y(n_2471)
);

INVx5_ASAP7_75t_L g2472 ( 
.A(n_2157),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2089),
.Y(n_2473)
);

BUFx3_ASAP7_75t_L g2474 ( 
.A(n_2158),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2089),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2080),
.Y(n_2476)
);

OAI21x1_ASAP7_75t_L g2477 ( 
.A1(n_2156),
.A2(n_1765),
.B(n_1725),
.Y(n_2477)
);

BUFx12f_ASAP7_75t_L g2478 ( 
.A(n_2067),
.Y(n_2478)
);

INVx3_ASAP7_75t_L g2479 ( 
.A(n_2081),
.Y(n_2479)
);

AOI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2135),
.A2(n_1341),
.B1(n_1342),
.B2(n_1339),
.Y(n_2480)
);

OA21x2_ASAP7_75t_L g2481 ( 
.A1(n_2065),
.A2(n_1814),
.B(n_1807),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2089),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_2205),
.B(n_1855),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2205),
.B(n_1858),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2089),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2089),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2089),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2089),
.Y(n_2488)
);

INVxp67_ASAP7_75t_L g2489 ( 
.A(n_2069),
.Y(n_2489)
);

OAI22x1_ASAP7_75t_SL g2490 ( 
.A1(n_2135),
.A2(n_1676),
.B1(n_1738),
.B2(n_1690),
.Y(n_2490)
);

BUFx6f_ASAP7_75t_L g2491 ( 
.A(n_2089),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2185),
.B(n_1869),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2094),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2080),
.B(n_1893),
.Y(n_2494)
);

OAI22x1_ASAP7_75t_L g2495 ( 
.A1(n_2134),
.A2(n_1823),
.B1(n_1917),
.B2(n_1655),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2089),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2089),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2205),
.B(n_1908),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2221),
.B(n_1455),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2070),
.Y(n_2500)
);

BUFx3_ASAP7_75t_L g2501 ( 
.A(n_2158),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2135),
.A2(n_1344),
.B1(n_1345),
.B2(n_1343),
.Y(n_2502)
);

BUFx12f_ASAP7_75t_L g2503 ( 
.A(n_2067),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2089),
.Y(n_2504)
);

AOI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2135),
.A2(n_1355),
.B1(n_1356),
.B2(n_1350),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2089),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2089),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2089),
.Y(n_2508)
);

INVx3_ASAP7_75t_L g2509 ( 
.A(n_2081),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2089),
.Y(n_2510)
);

INVx3_ASAP7_75t_L g2511 ( 
.A(n_2081),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2080),
.B(n_1906),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2205),
.B(n_1308),
.Y(n_2513)
);

BUFx6f_ASAP7_75t_L g2514 ( 
.A(n_2089),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2185),
.B(n_1933),
.Y(n_2515)
);

HB1xp67_ASAP7_75t_L g2516 ( 
.A(n_2094),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2089),
.Y(n_2517)
);

INVx3_ASAP7_75t_L g2518 ( 
.A(n_2081),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2069),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2135),
.A2(n_1363),
.B1(n_1370),
.B2(n_1360),
.Y(n_2520)
);

CKINVDCx6p67_ASAP7_75t_R g2521 ( 
.A(n_2221),
.Y(n_2521)
);

AND2x4_ASAP7_75t_L g2522 ( 
.A(n_2205),
.B(n_1954),
.Y(n_2522)
);

INVx5_ASAP7_75t_L g2523 ( 
.A(n_2157),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2089),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2089),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2089),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2089),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2205),
.B(n_1316),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2205),
.B(n_1329),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2205),
.B(n_1966),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2080),
.B(n_1985),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2089),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2089),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2089),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2205),
.B(n_1394),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2080),
.B(n_2009),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2089),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2089),
.Y(n_2538)
);

BUFx12f_ASAP7_75t_L g2539 ( 
.A(n_2067),
.Y(n_2539)
);

OA21x2_ASAP7_75t_L g2540 ( 
.A1(n_2065),
.A2(n_2033),
.B(n_2022),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2089),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2089),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_L g2543 ( 
.A(n_2185),
.B(n_2040),
.Y(n_2543)
);

AOI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_2135),
.A2(n_1377),
.B1(n_1388),
.B2(n_1374),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2081),
.Y(n_2545)
);

INVxp67_ASAP7_75t_L g2546 ( 
.A(n_2069),
.Y(n_2546)
);

OA21x2_ASAP7_75t_L g2547 ( 
.A1(n_2065),
.A2(n_2051),
.B(n_2045),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2081),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2135),
.A2(n_1390),
.B1(n_1392),
.B2(n_1389),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2185),
.B(n_1366),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2205),
.B(n_1520),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2080),
.B(n_1368),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2089),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2089),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2089),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_2089),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2351),
.Y(n_2557)
);

CKINVDCx20_ASAP7_75t_R g2558 ( 
.A(n_2500),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2369),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_2254),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2372),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2376),
.Y(n_2562)
);

BUFx10_ASAP7_75t_L g2563 ( 
.A(n_2401),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2377),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2253),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2256),
.Y(n_2566)
);

AND2x4_ASAP7_75t_L g2567 ( 
.A(n_2392),
.B(n_1566),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2399),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2408),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2381),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2382),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2425),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2417),
.B(n_1731),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2320),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2375),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2358),
.B(n_1455),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2327),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2330),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2268),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2447),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2448),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2364),
.B(n_1989),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2340),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2471),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2285),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2422),
.B(n_1756),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2344),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2353),
.Y(n_2588)
);

AND2x6_ASAP7_75t_L g2589 ( 
.A(n_2362),
.B(n_1435),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2333),
.B(n_1369),
.Y(n_2590)
);

CKINVDCx20_ASAP7_75t_R g2591 ( 
.A(n_2373),
.Y(n_2591)
);

CKINVDCx16_ASAP7_75t_R g2592 ( 
.A(n_2247),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2316),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2331),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2335),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2485),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_L g2597 ( 
.A(n_2487),
.Y(n_2597)
);

CKINVDCx20_ASAP7_75t_R g2598 ( 
.A(n_2329),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2398),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2413),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_2418),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2363),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_2426),
.Y(n_2603)
);

CKINVDCx20_ASAP7_75t_R g2604 ( 
.A(n_2521),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2367),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2325),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2488),
.Y(n_2607)
);

BUFx2_ASAP7_75t_L g2608 ( 
.A(n_2347),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2328),
.Y(n_2609)
);

NAND2x1_ASAP7_75t_L g2610 ( 
.A(n_2229),
.B(n_1435),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2491),
.Y(n_2611)
);

BUFx6f_ASAP7_75t_L g2612 ( 
.A(n_2504),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2338),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2384),
.Y(n_2614)
);

BUFx2_ASAP7_75t_L g2615 ( 
.A(n_2368),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2397),
.Y(n_2616)
);

INVx4_ASAP7_75t_L g2617 ( 
.A(n_2282),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2318),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_2454),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2378),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2507),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2239),
.B(n_1371),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2336),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2366),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2255),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2342),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2343),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2444),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2346),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2293),
.B(n_1375),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2232),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2299),
.B(n_1815),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2460),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2284),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2467),
.Y(n_2635)
);

INVxp67_ASAP7_75t_SL g2636 ( 
.A(n_2317),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2508),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2514),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2355),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2304),
.B(n_1380),
.Y(n_2640)
);

BUFx6f_ASAP7_75t_L g2641 ( 
.A(n_2517),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2478),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2463),
.B(n_1879),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2371),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2394),
.Y(n_2645)
);

INVx4_ASAP7_75t_L g2646 ( 
.A(n_2321),
.Y(n_2646)
);

BUFx2_ASAP7_75t_L g2647 ( 
.A(n_2240),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2474),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2264),
.A2(n_1776),
.B1(n_1816),
.B2(n_1803),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2277),
.B(n_1400),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2525),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2519),
.B(n_2043),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2501),
.Y(n_2653)
);

CKINVDCx6p67_ASAP7_75t_R g2654 ( 
.A(n_2235),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2503),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2348),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2352),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2526),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2555),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_L g2660 ( 
.A(n_2556),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2539),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2361),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2389),
.B(n_1521),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_L g2664 ( 
.A(n_2270),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2230),
.Y(n_2665)
);

CKINVDCx20_ASAP7_75t_R g2666 ( 
.A(n_2441),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2416),
.B(n_1399),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2379),
.Y(n_2668)
);

CKINVDCx20_ASAP7_75t_R g2669 ( 
.A(n_2275),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2283),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2326),
.Y(n_2671)
);

OR2x6_ASAP7_75t_L g2672 ( 
.A(n_2279),
.B(n_1564),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2431),
.B(n_1403),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_2345),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2432),
.B(n_1401),
.Y(n_2675)
);

CKINVDCx20_ASAP7_75t_R g2676 ( 
.A(n_2400),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2380),
.Y(n_2677)
);

HB1xp67_ASAP7_75t_L g2678 ( 
.A(n_2231),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2387),
.Y(n_2679)
);

HB1xp67_ASAP7_75t_L g2680 ( 
.A(n_2434),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2236),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2272),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2493),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_2267),
.Y(n_2684)
);

CKINVDCx20_ASAP7_75t_R g2685 ( 
.A(n_2516),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2324),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2259),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_R g2688 ( 
.A(n_2334),
.B(n_1405),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2402),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2357),
.B(n_1521),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2237),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2337),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2414),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2409),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2440),
.Y(n_2695)
);

CKINVDCx8_ASAP7_75t_R g2696 ( 
.A(n_2243),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2476),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2429),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2437),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2465),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2238),
.Y(n_2701)
);

BUFx3_ASAP7_75t_L g2702 ( 
.A(n_2385),
.Y(n_2702)
);

BUFx10_ASAP7_75t_L g2703 ( 
.A(n_2242),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2411),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2479),
.Y(n_2705)
);

BUFx3_ASAP7_75t_L g2706 ( 
.A(n_2386),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2509),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2412),
.Y(n_2708)
);

HB1xp67_ASAP7_75t_L g2709 ( 
.A(n_2234),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2245),
.Y(n_2710)
);

BUFx2_ASAP7_75t_L g2711 ( 
.A(n_2250),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2511),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2550),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2419),
.Y(n_2714)
);

OA21x2_ASAP7_75t_L g2715 ( 
.A1(n_2233),
.A2(n_1414),
.B(n_1407),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2435),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_2388),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2433),
.B(n_1416),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2449),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2457),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2518),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2486),
.Y(n_2722)
);

INVx1_ASAP7_75t_SL g2723 ( 
.A(n_2356),
.Y(n_2723)
);

CKINVDCx20_ASAP7_75t_R g2724 ( 
.A(n_2252),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_R g2725 ( 
.A(n_2251),
.B(n_2442),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2472),
.B(n_1428),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2545),
.Y(n_2727)
);

OA21x2_ASAP7_75t_L g2728 ( 
.A1(n_2262),
.A2(n_1468),
.B(n_1456),
.Y(n_2728)
);

HB1xp67_ASAP7_75t_L g2729 ( 
.A(n_2360),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2286),
.Y(n_2730)
);

INVx5_ASAP7_75t_L g2731 ( 
.A(n_2288),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2548),
.Y(n_2732)
);

CKINVDCx20_ASAP7_75t_R g2733 ( 
.A(n_2552),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2489),
.Y(n_2734)
);

OA21x2_ASAP7_75t_L g2735 ( 
.A1(n_2307),
.A2(n_1485),
.B(n_1473),
.Y(n_2735)
);

CKINVDCx16_ASAP7_75t_R g2736 ( 
.A(n_2246),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2374),
.Y(n_2737)
);

HB1xp67_ASAP7_75t_L g2738 ( 
.A(n_2428),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2301),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2523),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2496),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2311),
.Y(n_2742)
);

INVx6_ASAP7_75t_L g2743 ( 
.A(n_2294),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2506),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2248),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2461),
.B(n_1493),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2430),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2510),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2403),
.B(n_1427),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2261),
.Y(n_2750)
);

AND2x4_ASAP7_75t_L g2751 ( 
.A(n_2404),
.B(n_1429),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2527),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2468),
.B(n_1496),
.Y(n_2753)
);

BUFx8_ASAP7_75t_L g2754 ( 
.A(n_2249),
.Y(n_2754)
);

BUFx2_ASAP7_75t_L g2755 ( 
.A(n_2546),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2494),
.B(n_1404),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2280),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2339),
.B(n_1649),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_SL g2759 ( 
.A(n_2492),
.B(n_2515),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2498),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2410),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2289),
.Y(n_2762)
);

BUFx10_ASAP7_75t_L g2763 ( 
.A(n_2543),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2405),
.B(n_1432),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2534),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2271),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2257),
.B(n_1649),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2291),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2393),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2263),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2537),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2298),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2292),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2513),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2538),
.Y(n_2775)
);

INVxp67_ASAP7_75t_L g2776 ( 
.A(n_2528),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2295),
.Y(n_2777)
);

CKINVDCx20_ASAP7_75t_R g2778 ( 
.A(n_2499),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2541),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2300),
.Y(n_2780)
);

INVx6_ASAP7_75t_L g2781 ( 
.A(n_2365),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2512),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_2341),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2302),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_2531),
.Y(n_2785)
);

CKINVDCx20_ASAP7_75t_R g2786 ( 
.A(n_2281),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2309),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2554),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2265),
.Y(n_2789)
);

OA21x2_ASAP7_75t_L g2790 ( 
.A1(n_2395),
.A2(n_1513),
.B(n_1510),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2266),
.B(n_2529),
.Y(n_2791)
);

NAND2xp33_ASAP7_75t_R g2792 ( 
.A(n_2350),
.B(n_1408),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_SL g2793 ( 
.A(n_2273),
.B(n_1862),
.Y(n_2793)
);

BUFx2_ASAP7_75t_L g2794 ( 
.A(n_2396),
.Y(n_2794)
);

BUFx8_ASAP7_75t_L g2795 ( 
.A(n_2396),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_SL g2796 ( 
.A(n_2438),
.B(n_1881),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2536),
.B(n_1514),
.Y(n_2797)
);

CKINVDCx5p33_ASAP7_75t_R g2798 ( 
.A(n_2520),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2319),
.B(n_1519),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2535),
.B(n_1672),
.Y(n_2800)
);

XOR2xp5_ASAP7_75t_L g2801 ( 
.A(n_2443),
.B(n_1523),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2438),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2354),
.B(n_1529),
.Y(n_2803)
);

OA21x2_ASAP7_75t_L g2804 ( 
.A1(n_2407),
.A2(n_1539),
.B(n_1532),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2296),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2455),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2306),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2323),
.B(n_1545),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2310),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2269),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2480),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2258),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2391),
.B(n_1553),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2415),
.B(n_1557),
.Y(n_2814)
);

HB1xp67_ASAP7_75t_L g2815 ( 
.A(n_2551),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2260),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2423),
.B(n_1568),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2502),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2410),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2427),
.B(n_1571),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2278),
.Y(n_2821)
);

CKINVDCx20_ASAP7_75t_R g2822 ( 
.A(n_2505),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2274),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2544),
.B(n_1586),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2276),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2332),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2549),
.Y(n_2827)
);

NAND2xp33_ASAP7_75t_SL g2828 ( 
.A(n_2495),
.B(n_1882),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_2349),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2359),
.Y(n_2830)
);

CKINVDCx5p33_ASAP7_75t_R g2831 ( 
.A(n_2312),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2287),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_2322),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2313),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2314),
.Y(n_2835)
);

INVx3_ASAP7_75t_L g2836 ( 
.A(n_2436),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2477),
.Y(n_2837)
);

BUFx6f_ASAP7_75t_L g2838 ( 
.A(n_2436),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2450),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2490),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2459),
.B(n_2470),
.Y(n_2841)
);

BUFx2_ASAP7_75t_L g2842 ( 
.A(n_2483),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2290),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2484),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2303),
.Y(n_2845)
);

OAI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2522),
.A2(n_1412),
.B1(n_1413),
.B2(n_1411),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2530),
.B(n_1587),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2305),
.Y(n_2848)
);

OA21x2_ASAP7_75t_L g2849 ( 
.A1(n_2383),
.A2(n_2315),
.B(n_2308),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2241),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2244),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2406),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2420),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2297),
.Y(n_2854)
);

INVxp67_ASAP7_75t_L g2855 ( 
.A(n_2466),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2421),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2424),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2445),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2452),
.B(n_1417),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_2453),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2456),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2439),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2458),
.B(n_2462),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2469),
.Y(n_2864)
);

HB1xp67_ASAP7_75t_L g2865 ( 
.A(n_2370),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2390),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2473),
.Y(n_2867)
);

NAND2xp33_ASAP7_75t_R g2868 ( 
.A(n_2446),
.B(n_1419),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2475),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2482),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2560),
.Y(n_2871)
);

AND3x2_ASAP7_75t_L g2872 ( 
.A(n_2759),
.B(n_1282),
.C(n_1274),
.Y(n_2872)
);

BUFx2_ASAP7_75t_L g2873 ( 
.A(n_2669),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2863),
.Y(n_2874)
);

HB1xp67_ASAP7_75t_L g2875 ( 
.A(n_2709),
.Y(n_2875)
);

OR2x2_ASAP7_75t_SL g2876 ( 
.A(n_2592),
.B(n_1636),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2782),
.B(n_1596),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2558),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2557),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2559),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2665),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2691),
.Y(n_2882)
);

INVx3_ASAP7_75t_L g2883 ( 
.A(n_2807),
.Y(n_2883)
);

BUFx6f_ASAP7_75t_L g2884 ( 
.A(n_2560),
.Y(n_2884)
);

BUFx3_ASAP7_75t_L g2885 ( 
.A(n_2664),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2561),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2785),
.B(n_2451),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2750),
.B(n_2464),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2562),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2766),
.B(n_2481),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2865),
.A2(n_2540),
.B1(n_2547),
.B2(n_1702),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2701),
.Y(n_2892)
);

BUFx6f_ASAP7_75t_L g2893 ( 
.A(n_2568),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2704),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2564),
.Y(n_2895)
);

INVx3_ASAP7_75t_L g2896 ( 
.A(n_2568),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2570),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2580),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2768),
.B(n_1609),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2667),
.B(n_1621),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2675),
.B(n_1629),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2708),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2791),
.B(n_2713),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2800),
.B(n_2576),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2571),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2756),
.B(n_1632),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2663),
.B(n_2497),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2664),
.Y(n_2908)
);

INVx5_ASAP7_75t_L g2909 ( 
.A(n_2563),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2714),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2774),
.B(n_1634),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2776),
.B(n_1421),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2763),
.B(n_1422),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2866),
.A2(n_1702),
.B1(n_1378),
.B2(n_1418),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2632),
.B(n_1660),
.Y(n_2915)
);

INVxp33_ASAP7_75t_L g2916 ( 
.A(n_2582),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2870),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2710),
.Y(n_2918)
);

BUFx6f_ASAP7_75t_L g2919 ( 
.A(n_2580),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2793),
.B(n_1670),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2723),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_2739),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2716),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2719),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2596),
.Y(n_2925)
);

NAND3xp33_ASAP7_75t_L g2926 ( 
.A(n_2590),
.B(n_1424),
.C(n_1423),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2745),
.Y(n_2927)
);

INVx4_ASAP7_75t_L g2928 ( 
.A(n_2739),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2673),
.B(n_1425),
.Y(n_2929)
);

NAND2xp33_ASAP7_75t_SL g2930 ( 
.A(n_2688),
.B(n_1907),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2579),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2606),
.A2(n_1702),
.B1(n_1448),
.B2(n_1499),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2622),
.A2(n_1679),
.B1(n_1680),
.B2(n_1675),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2757),
.Y(n_2934)
);

NAND2xp33_ASAP7_75t_L g2935 ( 
.A(n_2589),
.B(n_1681),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2762),
.Y(n_2936)
);

BUFx2_ASAP7_75t_L g2937 ( 
.A(n_2674),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2803),
.B(n_1688),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2596),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2746),
.B(n_1693),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2773),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2720),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2753),
.B(n_1694),
.Y(n_2943)
);

BUFx3_ASAP7_75t_L g2944 ( 
.A(n_2742),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2585),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2777),
.Y(n_2946)
);

OAI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2796),
.A2(n_2833),
.B1(n_2831),
.B2(n_2806),
.Y(n_2947)
);

OR2x2_ASAP7_75t_L g2948 ( 
.A(n_2729),
.B(n_2524),
.Y(n_2948)
);

INVxp67_ASAP7_75t_L g2949 ( 
.A(n_2690),
.Y(n_2949)
);

BUFx2_ASAP7_75t_L g2950 ( 
.A(n_2676),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2780),
.Y(n_2951)
);

BUFx3_ASAP7_75t_L g2952 ( 
.A(n_2742),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2784),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2787),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2809),
.Y(n_2955)
);

OAI21xp33_ASAP7_75t_SL g2956 ( 
.A1(n_2636),
.A2(n_1438),
.B(n_1434),
.Y(n_2956)
);

BUFx8_ASAP7_75t_SL g2957 ( 
.A(n_2616),
.Y(n_2957)
);

HB1xp67_ASAP7_75t_L g2958 ( 
.A(n_2680),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2797),
.B(n_1433),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_SL g2960 ( 
.A1(n_2649),
.A2(n_2805),
.B1(n_2818),
.B2(n_2811),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2767),
.B(n_1710),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2722),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2741),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2630),
.B(n_1714),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2744),
.Y(n_2965)
);

AND2x2_ASAP7_75t_SL g2966 ( 
.A(n_2794),
.B(n_2647),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2748),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2640),
.B(n_1436),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2752),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2765),
.Y(n_2970)
);

INVxp67_ASAP7_75t_SL g2971 ( 
.A(n_2609),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2597),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2771),
.Y(n_2973)
);

INVx3_ASAP7_75t_L g2974 ( 
.A(n_2597),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2775),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2613),
.B(n_1739),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2779),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2589),
.A2(n_1702),
.B1(n_1501),
.B2(n_1559),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2788),
.Y(n_2979)
);

BUFx10_ASAP7_75t_L g2980 ( 
.A(n_2575),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2612),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2758),
.B(n_1753),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2656),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2607),
.B(n_2532),
.Y(n_2984)
);

AND3x2_ASAP7_75t_L g2985 ( 
.A(n_2711),
.B(n_1570),
.C(n_1294),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2618),
.B(n_1763),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2769),
.B(n_1437),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2789),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2623),
.B(n_1781),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2684),
.B(n_1784),
.Y(n_2990)
);

INVxp67_ASAP7_75t_L g2991 ( 
.A(n_2792),
.Y(n_2991)
);

BUFx2_ASAP7_75t_L g2992 ( 
.A(n_2685),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2626),
.B(n_1790),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2612),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2810),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2686),
.B(n_1795),
.Y(n_2996)
);

AND2x4_ASAP7_75t_L g2997 ( 
.A(n_2621),
.B(n_2533),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2657),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2627),
.B(n_1797),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2662),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2823),
.Y(n_3001)
);

INVx4_ASAP7_75t_L g3002 ( 
.A(n_2641),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2629),
.B(n_1800),
.Y(n_3003)
);

XOR2xp5_ASAP7_75t_L g3004 ( 
.A(n_2591),
.B(n_2614),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2815),
.B(n_2542),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2668),
.Y(n_3006)
);

AND2x6_ASAP7_75t_L g3007 ( 
.A(n_2837),
.B(n_1462),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2849),
.B(n_1817),
.Y(n_3008)
);

OR2x2_ASAP7_75t_L g3009 ( 
.A(n_2683),
.B(n_2553),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2677),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2738),
.B(n_1672),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2692),
.B(n_1818),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2679),
.Y(n_3013)
);

NAND3xp33_ASAP7_75t_L g3014 ( 
.A(n_2678),
.B(n_1443),
.C(n_1439),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2829),
.B(n_1444),
.Y(n_3015)
);

INVx2_ASAP7_75t_SL g3016 ( 
.A(n_2702),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2851),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2650),
.B(n_1830),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_2706),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2825),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2858),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2747),
.B(n_1747),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2832),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2850),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_L g3025 ( 
.A(n_2641),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2852),
.Y(n_3026)
);

AOI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2868),
.A2(n_1849),
.B1(n_1857),
.B2(n_1847),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2843),
.Y(n_3028)
);

INVx5_ASAP7_75t_L g3029 ( 
.A(n_2819),
.Y(n_3029)
);

NAND2xp33_ASAP7_75t_L g3030 ( 
.A(n_2589),
.B(n_2798),
.Y(n_3030)
);

BUFx3_ASAP7_75t_L g3031 ( 
.A(n_2658),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2841),
.A2(n_1874),
.B1(n_1889),
.B2(n_1872),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2760),
.B(n_1445),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2813),
.B(n_1901),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2848),
.Y(n_3035)
);

INVx4_ASAP7_75t_SL g3036 ( 
.A(n_2743),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2853),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2734),
.B(n_1747),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2808),
.B(n_1902),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_L g3040 ( 
.A(n_2827),
.B(n_1446),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2856),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_2717),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2857),
.Y(n_3043)
);

INVx2_ASAP7_75t_SL g3044 ( 
.A(n_2567),
.Y(n_3044)
);

INVx2_ASAP7_75t_SL g3045 ( 
.A(n_2573),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2658),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2864),
.Y(n_3047)
);

BUFx2_ASAP7_75t_L g3048 ( 
.A(n_2672),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2755),
.B(n_1447),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2694),
.B(n_1449),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2695),
.B(n_1911),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_SL g3052 ( 
.A(n_2593),
.B(n_1929),
.Y(n_3052)
);

INVx3_ASAP7_75t_L g3053 ( 
.A(n_2660),
.Y(n_3053)
);

INVx1_ASAP7_75t_SL g3054 ( 
.A(n_2615),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2867),
.Y(n_3055)
);

BUFx2_ASAP7_75t_L g3056 ( 
.A(n_2672),
.Y(n_3056)
);

BUFx10_ASAP7_75t_L g3057 ( 
.A(n_2625),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_2824),
.A2(n_1640),
.B1(n_1743),
.B2(n_1606),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2812),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_SL g3060 ( 
.A(n_2697),
.B(n_1913),
.Y(n_3060)
);

NAND2xp33_ASAP7_75t_SL g3061 ( 
.A(n_2786),
.B(n_1944),
.Y(n_3061)
);

AND2x4_ASAP7_75t_L g3062 ( 
.A(n_2569),
.B(n_2572),
.Y(n_3062)
);

AND2x6_ASAP7_75t_L g3063 ( 
.A(n_2631),
.B(n_1462),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2816),
.Y(n_3064)
);

OR2x6_ASAP7_75t_L g3065 ( 
.A(n_2781),
.B(n_1442),
.Y(n_3065)
);

BUFx3_ASAP7_75t_L g3066 ( 
.A(n_2660),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2845),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2565),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2860),
.B(n_1914),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2861),
.B(n_1920),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2681),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2687),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2689),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2693),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2733),
.B(n_1452),
.Y(n_3075)
);

BUFx2_ASAP7_75t_L g3076 ( 
.A(n_2670),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2698),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_2671),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2699),
.Y(n_3079)
);

BUFx6f_ASAP7_75t_L g3080 ( 
.A(n_2819),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2799),
.B(n_1921),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2700),
.Y(n_3082)
);

AND3x2_ASAP7_75t_L g3083 ( 
.A(n_2608),
.B(n_1766),
.C(n_1754),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2705),
.Y(n_3084)
);

NOR3xp33_ASAP7_75t_L g3085 ( 
.A(n_2828),
.B(n_2846),
.C(n_2842),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2707),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2839),
.B(n_1782),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2712),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2855),
.B(n_1923),
.Y(n_3089)
);

BUFx4f_ASAP7_75t_L g3090 ( 
.A(n_2654),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2721),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2869),
.B(n_1931),
.Y(n_3092)
);

BUFx8_ASAP7_75t_SL g3093 ( 
.A(n_2598),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2727),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2732),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_2682),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2749),
.A2(n_1821),
.B1(n_1831),
.B2(n_1810),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2834),
.Y(n_3098)
);

AOI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2854),
.A2(n_1961),
.B1(n_1986),
.B2(n_1934),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2835),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2826),
.Y(n_3101)
);

INVx3_ASAP7_75t_L g3102 ( 
.A(n_2566),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2586),
.B(n_1782),
.Y(n_3103)
);

INVx3_ASAP7_75t_L g3104 ( 
.A(n_2581),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_2584),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2830),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_2643),
.B(n_1454),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2611),
.Y(n_3108)
);

INVx2_ASAP7_75t_SL g3109 ( 
.A(n_2652),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2634),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2637),
.Y(n_3111)
);

BUFx6f_ASAP7_75t_L g3112 ( 
.A(n_2838),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2879),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2904),
.B(n_2594),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_2921),
.B(n_2916),
.Y(n_3115)
);

OAI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2887),
.A2(n_2822),
.B1(n_2817),
.B2(n_2820),
.Y(n_3116)
);

INVx2_ASAP7_75t_SL g3117 ( 
.A(n_2948),
.Y(n_3117)
);

INVx2_ASAP7_75t_SL g3118 ( 
.A(n_3009),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2880),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2991),
.B(n_2595),
.Y(n_3120)
);

AND2x2_ASAP7_75t_SL g3121 ( 
.A(n_3052),
.B(n_2736),
.Y(n_3121)
);

AO22x2_ASAP7_75t_L g3122 ( 
.A1(n_3085),
.A2(n_2801),
.B1(n_2764),
.B2(n_2751),
.Y(n_3122)
);

BUFx2_ASAP7_75t_L g3123 ( 
.A(n_2958),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2886),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2949),
.B(n_2599),
.Y(n_3125)
);

INVxp67_ASAP7_75t_SL g3126 ( 
.A(n_2893),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2968),
.B(n_2737),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2889),
.Y(n_3128)
);

INVxp67_ASAP7_75t_L g3129 ( 
.A(n_3038),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2929),
.B(n_2959),
.Y(n_3130)
);

HB1xp67_ASAP7_75t_L g3131 ( 
.A(n_2875),
.Y(n_3131)
);

AND2x4_ASAP7_75t_L g3132 ( 
.A(n_2909),
.B(n_2639),
.Y(n_3132)
);

BUFx4f_ASAP7_75t_L g3133 ( 
.A(n_3080),
.Y(n_3133)
);

INVx4_ASAP7_75t_L g3134 ( 
.A(n_2909),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2982),
.B(n_2600),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2895),
.Y(n_3136)
);

BUFx4f_ASAP7_75t_L g3137 ( 
.A(n_3080),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2881),
.Y(n_3138)
);

OR2x2_ASAP7_75t_SL g3139 ( 
.A(n_3042),
.B(n_2814),
.Y(n_3139)
);

NAND2x1p5_ASAP7_75t_L g3140 ( 
.A(n_2883),
.B(n_2731),
.Y(n_3140)
);

INVxp67_ASAP7_75t_L g3141 ( 
.A(n_3049),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_3112),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2882),
.Y(n_3143)
);

AOI22xp33_ASAP7_75t_L g3144 ( 
.A1(n_2888),
.A2(n_2802),
.B1(n_2610),
.B2(n_2645),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2897),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2905),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_2931),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2892),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2874),
.B(n_2601),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2927),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_R g3151 ( 
.A(n_2945),
.B(n_2603),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2894),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2934),
.Y(n_3153)
);

BUFx6f_ASAP7_75t_L g3154 ( 
.A(n_3112),
.Y(n_3154)
);

AND2x2_ASAP7_75t_SL g3155 ( 
.A(n_3076),
.B(n_2646),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2902),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2910),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2936),
.Y(n_3158)
);

INVx4_ASAP7_75t_L g3159 ( 
.A(n_3029),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_2890),
.A2(n_2648),
.B1(n_2653),
.B2(n_2644),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2941),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2923),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_3015),
.B(n_2847),
.Y(n_3163)
);

INVxp67_ASAP7_75t_L g3164 ( 
.A(n_3011),
.Y(n_3164)
);

BUFx2_ASAP7_75t_L g3165 ( 
.A(n_2873),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_3040),
.B(n_2703),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2924),
.Y(n_3167)
);

INVx5_ASAP7_75t_L g3168 ( 
.A(n_2957),
.Y(n_3168)
);

OAI22xp5_ASAP7_75t_SL g3169 ( 
.A1(n_2960),
.A2(n_2619),
.B1(n_2783),
.B2(n_2778),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_2903),
.B(n_2844),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2900),
.B(n_2821),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2871),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_SL g3173 ( 
.A(n_3078),
.B(n_2628),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2946),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2951),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_L g3176 ( 
.A1(n_2953),
.A2(n_2859),
.B1(n_2804),
.B2(n_1462),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2901),
.B(n_2725),
.Y(n_3177)
);

AND2x4_ASAP7_75t_L g3178 ( 
.A(n_3036),
.B(n_2638),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2954),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2955),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2871),
.Y(n_3181)
);

BUFx2_ASAP7_75t_L g3182 ( 
.A(n_2937),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_2918),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3017),
.Y(n_3184)
);

NOR2x1p5_ASAP7_75t_L g3185 ( 
.A(n_2885),
.B(n_2633),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3021),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2962),
.Y(n_3187)
);

INVx3_ASAP7_75t_L g3188 ( 
.A(n_2893),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2942),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_3029),
.Y(n_3190)
);

NAND2x1p5_ASAP7_75t_L g3191 ( 
.A(n_2928),
.B(n_2731),
.Y(n_3191)
);

BUFx6f_ASAP7_75t_L g3192 ( 
.A(n_2884),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2907),
.B(n_2651),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_2950),
.Y(n_3194)
);

AO22x2_ASAP7_75t_L g3195 ( 
.A1(n_3004),
.A2(n_1466),
.B1(n_1467),
.B2(n_1461),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2947),
.B(n_2624),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_2884),
.Y(n_3197)
);

NAND3x1_ASAP7_75t_L g3198 ( 
.A(n_3075),
.B(n_2840),
.C(n_2666),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_L g3199 ( 
.A(n_2913),
.B(n_2718),
.Y(n_3199)
);

BUFx2_ASAP7_75t_L g3200 ( 
.A(n_2992),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2963),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2973),
.Y(n_3202)
);

BUFx3_ASAP7_75t_L g3203 ( 
.A(n_2898),
.Y(n_3203)
);

AO22x2_ASAP7_75t_L g3204 ( 
.A1(n_2917),
.A2(n_1500),
.B1(n_1504),
.B2(n_1475),
.Y(n_3204)
);

BUFx2_ASAP7_75t_L g3205 ( 
.A(n_2878),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2965),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_2906),
.B(n_2795),
.Y(n_3207)
);

HB1xp67_ASAP7_75t_L g3208 ( 
.A(n_3016),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3050),
.B(n_2659),
.Y(n_3209)
);

NAND3xp33_ASAP7_75t_L g3210 ( 
.A(n_3033),
.B(n_2726),
.C(n_2754),
.Y(n_3210)
);

BUFx2_ASAP7_75t_L g3211 ( 
.A(n_3019),
.Y(n_3211)
);

AND3x4_ASAP7_75t_L g3212 ( 
.A(n_2981),
.B(n_2772),
.C(n_2770),
.Y(n_3212)
);

AND2x6_ASAP7_75t_L g3213 ( 
.A(n_3110),
.B(n_1505),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2979),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_2898),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2919),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_2919),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_3096),
.B(n_2574),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2967),
.Y(n_3219)
);

NAND2x1p5_ASAP7_75t_L g3220 ( 
.A(n_3002),
.B(n_2730),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2969),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2988),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2987),
.B(n_2740),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2971),
.B(n_1987),
.Y(n_3224)
);

BUFx6f_ASAP7_75t_L g3225 ( 
.A(n_2972),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2972),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2940),
.B(n_1998),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2995),
.Y(n_3228)
);

BUFx3_ASAP7_75t_L g3229 ( 
.A(n_3025),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_2914),
.A2(n_1956),
.B1(n_1962),
.B2(n_1950),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2970),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2943),
.B(n_2000),
.Y(n_3232)
);

OAI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2891),
.A2(n_1996),
.B1(n_2006),
.B2(n_1978),
.Y(n_3233)
);

AND2x4_ASAP7_75t_L g3234 ( 
.A(n_2908),
.B(n_2577),
.Y(n_3234)
);

INVxp67_ASAP7_75t_L g3235 ( 
.A(n_3022),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_2877),
.B(n_2604),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_SL g3237 ( 
.A1(n_2876),
.A2(n_2021),
.B1(n_2024),
.B2(n_2019),
.Y(n_3237)
);

NAND3x1_ASAP7_75t_L g3238 ( 
.A(n_3099),
.B(n_1515),
.C(n_1507),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2975),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2899),
.B(n_2578),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_2912),
.B(n_3069),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2964),
.B(n_2002),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_3025),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3001),
.Y(n_3244)
);

BUFx2_ASAP7_75t_L g3245 ( 
.A(n_3046),
.Y(n_3245)
);

OAI22xp5_ASAP7_75t_SL g3246 ( 
.A1(n_2966),
.A2(n_2057),
.B1(n_2724),
.B2(n_2642),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2977),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2983),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3020),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3023),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_3046),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3028),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_2922),
.B(n_2583),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3035),
.Y(n_3254)
);

OAI22xp5_ASAP7_75t_SL g3255 ( 
.A1(n_3048),
.A2(n_2635),
.B1(n_2661),
.B2(n_2655),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_2944),
.Y(n_3256)
);

INVx4_ASAP7_75t_L g3257 ( 
.A(n_2994),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2915),
.B(n_2696),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2938),
.B(n_2017),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_3031),
.Y(n_3260)
);

INVx5_ASAP7_75t_L g3261 ( 
.A(n_3093),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3081),
.B(n_2587),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_3066),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2998),
.Y(n_3264)
);

INVxp67_ASAP7_75t_L g3265 ( 
.A(n_3087),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3000),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3006),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3068),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_2952),
.B(n_2588),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3034),
.B(n_2025),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3045),
.B(n_2602),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_3130),
.B(n_2930),
.Y(n_3272)
);

OR2x6_ASAP7_75t_L g3273 ( 
.A(n_3123),
.B(n_3065),
.Y(n_3273)
);

INVx3_ASAP7_75t_L g3274 ( 
.A(n_3159),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_3171),
.A2(n_3008),
.B(n_3039),
.Y(n_3275)
);

NAND3xp33_ASAP7_75t_SL g3276 ( 
.A(n_3166),
.B(n_3027),
.C(n_3061),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3241),
.B(n_3018),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_L g3278 ( 
.A1(n_3113),
.A2(n_3124),
.B1(n_3128),
.B2(n_3119),
.Y(n_3278)
);

INVx1_ASAP7_75t_SL g3279 ( 
.A(n_3115),
.Y(n_3279)
);

INVx5_ASAP7_75t_L g3280 ( 
.A(n_3142),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3127),
.B(n_2872),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_3142),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3138),
.Y(n_3283)
);

AND2x6_ASAP7_75t_SL g3284 ( 
.A(n_3236),
.B(n_3065),
.Y(n_3284)
);

A2O1A1Ixp33_ASAP7_75t_SL g3285 ( 
.A1(n_3199),
.A2(n_3030),
.B(n_3107),
.C(n_3067),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3141),
.B(n_3010),
.Y(n_3286)
);

INVxp67_ASAP7_75t_L g3287 ( 
.A(n_3131),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_SL g3288 ( 
.A(n_3147),
.B(n_3057),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_3163),
.B(n_3070),
.Y(n_3289)
);

BUFx2_ASAP7_75t_L g3290 ( 
.A(n_3165),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3143),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3177),
.B(n_3013),
.Y(n_3292)
);

INVxp67_ASAP7_75t_L g3293 ( 
.A(n_3117),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_SL g3294 ( 
.A(n_3116),
.B(n_3089),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_3151),
.B(n_2926),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3136),
.B(n_3024),
.Y(n_3296)
);

INVxp67_ASAP7_75t_L g3297 ( 
.A(n_3118),
.Y(n_3297)
);

A2O1A1Ixp33_ASAP7_75t_SL g3298 ( 
.A1(n_3240),
.A2(n_3064),
.B(n_3059),
.C(n_3071),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3145),
.B(n_3146),
.Y(n_3299)
);

AND2x4_ASAP7_75t_L g3300 ( 
.A(n_3256),
.B(n_3257),
.Y(n_3300)
);

INVx3_ASAP7_75t_L g3301 ( 
.A(n_3190),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_L g3302 ( 
.A(n_3120),
.B(n_3092),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3150),
.B(n_3153),
.Y(n_3303)
);

NOR2xp33_ASAP7_75t_L g3304 ( 
.A(n_3233),
.B(n_2990),
.Y(n_3304)
);

OR2x2_ASAP7_75t_L g3305 ( 
.A(n_3182),
.B(n_3005),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3158),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3161),
.B(n_3026),
.Y(n_3307)
);

NAND2x1p5_ASAP7_75t_L g3308 ( 
.A(n_3133),
.B(n_2896),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_3178),
.B(n_3109),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3174),
.Y(n_3310)
);

O2A1O1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_3164),
.A2(n_2920),
.B(n_2956),
.C(n_2961),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3175),
.B(n_3037),
.Y(n_3312)
);

AND2x6_ASAP7_75t_SL g3313 ( 
.A(n_3196),
.B(n_3103),
.Y(n_3313)
);

CKINVDCx5p33_ASAP7_75t_R g3314 ( 
.A(n_3261),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3148),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3179),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3125),
.B(n_2976),
.Y(n_3317)
);

INVxp67_ASAP7_75t_L g3318 ( 
.A(n_3183),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3155),
.B(n_2986),
.Y(n_3319)
);

BUFx6f_ASAP7_75t_L g3320 ( 
.A(n_3154),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3180),
.B(n_3047),
.Y(n_3321)
);

AND2x2_ASAP7_75t_L g3322 ( 
.A(n_3129),
.B(n_3044),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_3230),
.B(n_3235),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3184),
.Y(n_3324)
);

AND2x4_ASAP7_75t_L g3325 ( 
.A(n_3234),
.B(n_3253),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_3265),
.B(n_2996),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3186),
.B(n_3055),
.Y(n_3327)
);

NAND3xp33_ASAP7_75t_L g3328 ( 
.A(n_3223),
.B(n_3160),
.C(n_3014),
.Y(n_3328)
);

INVxp67_ASAP7_75t_L g3329 ( 
.A(n_3217),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_3209),
.B(n_2989),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3248),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3264),
.B(n_3041),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3266),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3267),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3152),
.Y(n_3335)
);

AOI21xp33_ASAP7_75t_L g3336 ( 
.A1(n_3224),
.A2(n_2911),
.B(n_3012),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_3245),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3156),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3187),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3157),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3227),
.B(n_3043),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_L g3342 ( 
.A1(n_3162),
.A2(n_3100),
.B1(n_3101),
.B2(n_3098),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_3269),
.B(n_2925),
.Y(n_3343)
);

NAND2xp33_ASAP7_75t_L g3344 ( 
.A(n_3144),
.B(n_3007),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3154),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_SL g3346 ( 
.A1(n_3121),
.A2(n_3056),
.B1(n_3106),
.B2(n_2980),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3193),
.B(n_3054),
.Y(n_3347)
);

AOI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_3135),
.A2(n_2933),
.B1(n_3060),
.B2(n_3051),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3206),
.Y(n_3349)
);

AOI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3114),
.A2(n_3032),
.B1(n_3073),
.B2(n_3072),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3219),
.Y(n_3351)
);

OR2x6_ASAP7_75t_L g3352 ( 
.A(n_3134),
.B(n_2939),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3167),
.A2(n_3088),
.B1(n_3091),
.B2(n_3079),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3189),
.Y(n_3354)
);

NOR2x1_ASAP7_75t_R g3355 ( 
.A(n_3168),
.B(n_2617),
.Y(n_3355)
);

CKINVDCx5p33_ASAP7_75t_R g3356 ( 
.A(n_3261),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_3194),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_3137),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_3218),
.B(n_3132),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3232),
.B(n_3094),
.Y(n_3360)
);

AND2x4_ASAP7_75t_L g3361 ( 
.A(n_3203),
.B(n_2974),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3173),
.B(n_2993),
.Y(n_3362)
);

NOR2x2_ASAP7_75t_L g3363 ( 
.A(n_3201),
.B(n_3202),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3242),
.B(n_3095),
.Y(n_3364)
);

CKINVDCx20_ASAP7_75t_R g3365 ( 
.A(n_3168),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3221),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_3215),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_3149),
.B(n_3074),
.Y(n_3368)
);

INVx1_ASAP7_75t_SL g3369 ( 
.A(n_3200),
.Y(n_3369)
);

O2A1O1Ixp33_ASAP7_75t_L g3370 ( 
.A1(n_3258),
.A2(n_2935),
.B(n_3003),
.C(n_2999),
.Y(n_3370)
);

INVxp67_ASAP7_75t_SL g3371 ( 
.A(n_3208),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_3211),
.B(n_3077),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3260),
.Y(n_3373)
);

AOI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3169),
.A2(n_3082),
.B1(n_3086),
.B2(n_3084),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3259),
.B(n_3058),
.Y(n_3375)
);

OAI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3231),
.A2(n_3111),
.B1(n_3108),
.B2(n_3105),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3204),
.B(n_3062),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3239),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3270),
.B(n_3097),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3205),
.B(n_3053),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_3214),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3247),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3222),
.B(n_3228),
.Y(n_3383)
);

OAI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3176),
.A2(n_2978),
.B1(n_2932),
.B2(n_3104),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_3172),
.Y(n_3385)
);

NOR2x2_ASAP7_75t_L g3386 ( 
.A(n_3244),
.B(n_1952),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3249),
.B(n_3007),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3172),
.B(n_2984),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3250),
.Y(n_3389)
);

AND2x6_ASAP7_75t_L g3390 ( 
.A(n_3181),
.B(n_3192),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3252),
.A2(n_3007),
.B1(n_2997),
.B2(n_1749),
.Y(n_3391)
);

AND2x2_ASAP7_75t_L g3392 ( 
.A(n_3126),
.B(n_3102),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3254),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3268),
.B(n_2605),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3262),
.B(n_2029),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3271),
.Y(n_3396)
);

AO22x1_ASAP7_75t_L g3397 ( 
.A1(n_3212),
.A2(n_2620),
.B1(n_1458),
.B2(n_1459),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3251),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_3170),
.B(n_3090),
.Y(n_3399)
);

CKINVDCx5p33_ASAP7_75t_R g3400 ( 
.A(n_3255),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3260),
.B(n_1457),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3188),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3216),
.Y(n_3403)
);

OR2x2_ASAP7_75t_L g3404 ( 
.A(n_3139),
.B(n_1460),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3306),
.Y(n_3405)
);

BUFx6f_ASAP7_75t_L g3406 ( 
.A(n_3320),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3277),
.B(n_3238),
.Y(n_3407)
);

INVxp33_ASAP7_75t_L g3408 ( 
.A(n_3347),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3323),
.B(n_3122),
.Y(n_3409)
);

BUFx6f_ASAP7_75t_L g3410 ( 
.A(n_3320),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3290),
.Y(n_3411)
);

INVx4_ASAP7_75t_L g3412 ( 
.A(n_3280),
.Y(n_3412)
);

AOI22xp33_ASAP7_75t_L g3413 ( 
.A1(n_3304),
.A2(n_3276),
.B1(n_3289),
.B2(n_3302),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3310),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3292),
.B(n_3263),
.Y(n_3415)
);

INVx3_ASAP7_75t_L g3416 ( 
.A(n_3300),
.Y(n_3416)
);

BUFx3_ASAP7_75t_L g3417 ( 
.A(n_3280),
.Y(n_3417)
);

BUFx3_ASAP7_75t_L g3418 ( 
.A(n_3358),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_3279),
.B(n_3246),
.Y(n_3419)
);

CKINVDCx20_ASAP7_75t_R g3420 ( 
.A(n_3365),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_3287),
.B(n_3237),
.Y(n_3421)
);

BUFx2_ASAP7_75t_L g3422 ( 
.A(n_3357),
.Y(n_3422)
);

INVx4_ASAP7_75t_L g3423 ( 
.A(n_3390),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3316),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_R g3425 ( 
.A(n_3288),
.B(n_3263),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3324),
.Y(n_3426)
);

INVx3_ASAP7_75t_L g3427 ( 
.A(n_3367),
.Y(n_3427)
);

INVx3_ASAP7_75t_L g3428 ( 
.A(n_3373),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3360),
.B(n_3140),
.Y(n_3429)
);

BUFx3_ASAP7_75t_L g3430 ( 
.A(n_3282),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3364),
.B(n_3181),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3281),
.B(n_3192),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_3305),
.B(n_3197),
.Y(n_3433)
);

NAND3xp33_ASAP7_75t_SL g3434 ( 
.A(n_3328),
.B(n_3207),
.C(n_3210),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3331),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3333),
.Y(n_3436)
);

NAND3xp33_ASAP7_75t_L g3437 ( 
.A(n_3272),
.B(n_2985),
.C(n_3083),
.Y(n_3437)
);

OR2x2_ASAP7_75t_L g3438 ( 
.A(n_3369),
.B(n_3229),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3334),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3286),
.B(n_3330),
.Y(n_3440)
);

AOI21xp33_ASAP7_75t_L g3441 ( 
.A1(n_3294),
.A2(n_3195),
.B(n_3198),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_3390),
.Y(n_3442)
);

BUFx4f_ASAP7_75t_L g3443 ( 
.A(n_3390),
.Y(n_3443)
);

CKINVDCx6p67_ASAP7_75t_R g3444 ( 
.A(n_3273),
.Y(n_3444)
);

AOI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3326),
.A2(n_3319),
.B1(n_3317),
.B2(n_3399),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_3325),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_R g3447 ( 
.A(n_3314),
.B(n_3197),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3339),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3299),
.B(n_3225),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_R g3450 ( 
.A(n_3356),
.B(n_3400),
.Y(n_3450)
);

NAND2x1_ASAP7_75t_L g3451 ( 
.A(n_3349),
.B(n_3225),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_L g3452 ( 
.A(n_3318),
.B(n_3226),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3303),
.B(n_3226),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3351),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3366),
.Y(n_3455)
);

BUFx3_ASAP7_75t_L g3456 ( 
.A(n_3359),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3293),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3361),
.Y(n_3458)
);

BUFx2_ASAP7_75t_L g3459 ( 
.A(n_3363),
.Y(n_3459)
);

CKINVDCx5p33_ASAP7_75t_R g3460 ( 
.A(n_3313),
.Y(n_3460)
);

INVx3_ASAP7_75t_L g3461 ( 
.A(n_3308),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3378),
.Y(n_3462)
);

INVx2_ASAP7_75t_SL g3463 ( 
.A(n_3385),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3343),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3377),
.A2(n_3185),
.B1(n_3213),
.B2(n_3063),
.Y(n_3465)
);

OR2x6_ASAP7_75t_L g3466 ( 
.A(n_3273),
.B(n_3243),
.Y(n_3466)
);

NOR3xp33_ASAP7_75t_SL g3467 ( 
.A(n_3295),
.B(n_1464),
.C(n_1463),
.Y(n_3467)
);

HB1xp67_ASAP7_75t_L g3468 ( 
.A(n_3297),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3382),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3278),
.B(n_3243),
.Y(n_3470)
);

INVx1_ASAP7_75t_SL g3471 ( 
.A(n_3386),
.Y(n_3471)
);

NOR3xp33_ASAP7_75t_SL g3472 ( 
.A(n_3362),
.B(n_1471),
.C(n_1469),
.Y(n_3472)
);

INVx3_ASAP7_75t_L g3473 ( 
.A(n_3274),
.Y(n_3473)
);

OAI221xp5_ASAP7_75t_L g3474 ( 
.A1(n_3346),
.A2(n_3220),
.B1(n_3191),
.B2(n_1527),
.C(n_1535),
.Y(n_3474)
);

CKINVDCx20_ASAP7_75t_R g3475 ( 
.A(n_3329),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3332),
.Y(n_3476)
);

INVx2_ASAP7_75t_SL g3477 ( 
.A(n_3345),
.Y(n_3477)
);

INVx2_ASAP7_75t_SL g3478 ( 
.A(n_3309),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_3284),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3341),
.B(n_3213),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3368),
.B(n_3213),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3283),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_3337),
.B(n_3398),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3374),
.B(n_1787),
.Y(n_3484)
);

AND2x2_ASAP7_75t_SL g3485 ( 
.A(n_3344),
.B(n_1505),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3296),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3275),
.A2(n_2728),
.B(n_2715),
.Y(n_3487)
);

INVxp67_ASAP7_75t_L g3488 ( 
.A(n_3401),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3307),
.Y(n_3489)
);

NOR3xp33_ASAP7_75t_SL g3490 ( 
.A(n_3388),
.B(n_1477),
.C(n_1476),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3312),
.Y(n_3491)
);

INVx2_ASAP7_75t_SL g3492 ( 
.A(n_3352),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3379),
.B(n_3063),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_3352),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3291),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_3322),
.Y(n_3496)
);

HB1xp67_ASAP7_75t_L g3497 ( 
.A(n_3371),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3321),
.Y(n_3498)
);

NOR3xp33_ASAP7_75t_SL g3499 ( 
.A(n_3380),
.B(n_1481),
.C(n_1480),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3396),
.B(n_3392),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3315),
.B(n_1787),
.Y(n_3501)
);

NAND2xp33_ASAP7_75t_R g3502 ( 
.A(n_3301),
.B(n_2735),
.Y(n_3502)
);

BUFx2_ASAP7_75t_L g3503 ( 
.A(n_3402),
.Y(n_3503)
);

HB1xp67_ASAP7_75t_L g3504 ( 
.A(n_3403),
.Y(n_3504)
);

CKINVDCx5p33_ASAP7_75t_R g3505 ( 
.A(n_3404),
.Y(n_3505)
);

INVx1_ASAP7_75t_SL g3506 ( 
.A(n_3372),
.Y(n_3506)
);

CKINVDCx8_ASAP7_75t_R g3507 ( 
.A(n_3355),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3348),
.A2(n_2037),
.B1(n_2046),
.B2(n_2031),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_3350),
.B(n_1793),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3413),
.B(n_3327),
.Y(n_3510)
);

AO31x2_ASAP7_75t_L g3511 ( 
.A1(n_3487),
.A2(n_3384),
.A3(n_3375),
.B(n_3387),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3486),
.B(n_3335),
.Y(n_3512)
);

AOI21xp33_ASAP7_75t_L g3513 ( 
.A1(n_3509),
.A2(n_3285),
.B(n_3311),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3485),
.A2(n_3370),
.B(n_3336),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3500),
.B(n_3408),
.Y(n_3515)
);

OAI22x1_ASAP7_75t_L g3516 ( 
.A1(n_3445),
.A2(n_3340),
.B1(n_3354),
.B2(n_3338),
.Y(n_3516)
);

BUFx2_ASAP7_75t_L g3517 ( 
.A(n_3475),
.Y(n_3517)
);

NAND3xp33_ASAP7_75t_SL g3518 ( 
.A(n_3488),
.B(n_3395),
.C(n_3353),
.Y(n_3518)
);

BUFx6f_ASAP7_75t_L g3519 ( 
.A(n_3417),
.Y(n_3519)
);

O2A1O1Ixp5_ASAP7_75t_L g3520 ( 
.A1(n_3484),
.A2(n_3441),
.B(n_3481),
.C(n_3407),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3489),
.A2(n_3298),
.B(n_2790),
.Y(n_3521)
);

AOI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_3491),
.A2(n_3391),
.B(n_3383),
.Y(n_3522)
);

BUFx3_ASAP7_75t_L g3523 ( 
.A(n_3418),
.Y(n_3523)
);

AND2x4_ASAP7_75t_L g3524 ( 
.A(n_3430),
.B(n_3381),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3429),
.B(n_3342),
.Y(n_3525)
);

A2O1A1Ixp33_ASAP7_75t_L g3526 ( 
.A1(n_3434),
.A2(n_3393),
.B(n_3389),
.C(n_3394),
.Y(n_3526)
);

OAI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3508),
.A2(n_3376),
.B(n_3063),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3498),
.B(n_3397),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3476),
.B(n_3440),
.Y(n_3529)
);

OAI21x1_ASAP7_75t_L g3530 ( 
.A1(n_3493),
.A2(n_1524),
.B(n_1522),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3424),
.Y(n_3531)
);

HB1xp67_ASAP7_75t_L g3532 ( 
.A(n_3457),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3480),
.A2(n_1749),
.B(n_1505),
.Y(n_3533)
);

AOI221xp5_ASAP7_75t_SL g3534 ( 
.A1(n_3474),
.A2(n_1546),
.B1(n_1547),
.B2(n_1538),
.C(n_1537),
.Y(n_3534)
);

AOI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3505),
.A2(n_2064),
.B1(n_1483),
.B2(n_1486),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3415),
.A2(n_1762),
.B(n_1749),
.Y(n_3536)
);

BUFx3_ASAP7_75t_L g3537 ( 
.A(n_3406),
.Y(n_3537)
);

OAI21x1_ASAP7_75t_L g3538 ( 
.A1(n_3405),
.A2(n_1561),
.B(n_1552),
.Y(n_3538)
);

NAND3xp33_ASAP7_75t_L g3539 ( 
.A(n_3467),
.B(n_1492),
.C(n_1482),
.Y(n_3539)
);

OAI21x1_ASAP7_75t_SL g3540 ( 
.A1(n_3470),
.A2(n_1963),
.B(n_1953),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3431),
.A2(n_1785),
.B(n_1762),
.Y(n_3541)
);

A2O1A1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3472),
.A2(n_1569),
.B(n_1574),
.C(n_1563),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3496),
.B(n_1494),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3435),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3506),
.B(n_1793),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3449),
.B(n_1498),
.Y(n_3546)
);

AOI21x1_ASAP7_75t_L g3547 ( 
.A1(n_3409),
.A2(n_1595),
.B(n_1588),
.Y(n_3547)
);

OAI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3414),
.A2(n_3436),
.B(n_3426),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3453),
.B(n_1503),
.Y(n_3549)
);

INVxp67_ASAP7_75t_L g3550 ( 
.A(n_3411),
.Y(n_3550)
);

AOI21xp33_ASAP7_75t_L g3551 ( 
.A1(n_3502),
.A2(n_1599),
.B(n_1597),
.Y(n_3551)
);

INVx3_ASAP7_75t_L g3552 ( 
.A(n_3412),
.Y(n_3552)
);

CKINVDCx5p33_ASAP7_75t_R g3553 ( 
.A(n_3425),
.Y(n_3553)
);

XNOR2xp5_ASAP7_75t_L g3554 ( 
.A(n_3420),
.B(n_1511),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_3450),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3446),
.B(n_1512),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3439),
.A2(n_1618),
.B(n_1612),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3421),
.B(n_1517),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3459),
.B(n_1518),
.Y(n_3559)
);

OAI22x1_ASAP7_75t_L g3560 ( 
.A1(n_3460),
.A2(n_1630),
.B1(n_1652),
.B2(n_1627),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3448),
.Y(n_3561)
);

BUFx6f_ASAP7_75t_L g3562 ( 
.A(n_3406),
.Y(n_3562)
);

AOI21xp5_ASAP7_75t_L g3563 ( 
.A1(n_3455),
.A2(n_1785),
.B(n_1762),
.Y(n_3563)
);

AOI21x1_ASAP7_75t_L g3564 ( 
.A1(n_3451),
.A2(n_1654),
.B(n_1653),
.Y(n_3564)
);

OAI21x1_ASAP7_75t_L g3565 ( 
.A1(n_3454),
.A2(n_1682),
.B(n_1664),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3462),
.A2(n_1928),
.B(n_1785),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3432),
.B(n_1525),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3416),
.B(n_1536),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3419),
.B(n_1544),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3501),
.B(n_1548),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3469),
.A2(n_2038),
.B(n_1928),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3482),
.A2(n_1697),
.B(n_1695),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3495),
.Y(n_3573)
);

BUFx2_ASAP7_75t_L g3574 ( 
.A(n_3422),
.Y(n_3574)
);

AO31x2_ASAP7_75t_L g3575 ( 
.A1(n_3503),
.A2(n_2023),
.A3(n_2050),
.B(n_2012),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3497),
.B(n_1549),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3468),
.B(n_3464),
.Y(n_3577)
);

OAI21x1_ASAP7_75t_L g3578 ( 
.A1(n_3433),
.A2(n_1723),
.B(n_1721),
.Y(n_3578)
);

OA21x2_ASAP7_75t_L g3579 ( 
.A1(n_3437),
.A2(n_1737),
.B(n_1735),
.Y(n_3579)
);

INVx3_ASAP7_75t_L g3580 ( 
.A(n_3427),
.Y(n_3580)
);

AOI21xp33_ASAP7_75t_L g3581 ( 
.A1(n_3504),
.A2(n_1750),
.B(n_1742),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3443),
.A2(n_3465),
.B(n_3466),
.Y(n_3582)
);

OAI21x1_ASAP7_75t_L g3583 ( 
.A1(n_3461),
.A2(n_1760),
.B(n_1758),
.Y(n_3583)
);

AOI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3466),
.A2(n_2038),
.B(n_1928),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3483),
.B(n_1550),
.Y(n_3585)
);

OAI21x1_ASAP7_75t_L g3586 ( 
.A1(n_3473),
.A2(n_1764),
.B(n_1761),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3463),
.Y(n_3587)
);

INVx1_ASAP7_75t_SL g3588 ( 
.A(n_3438),
.Y(n_3588)
);

O2A1O1Ixp5_ASAP7_75t_L g3589 ( 
.A1(n_3452),
.A2(n_1786),
.B(n_1788),
.C(n_1780),
.Y(n_3589)
);

OA21x2_ASAP7_75t_L g3590 ( 
.A1(n_3490),
.A2(n_1798),
.B(n_1792),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3478),
.B(n_3456),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3458),
.B(n_1554),
.Y(n_3592)
);

OAI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3499),
.A2(n_1808),
.B(n_1804),
.Y(n_3593)
);

HB1xp67_ASAP7_75t_L g3594 ( 
.A(n_3410),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3492),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3428),
.Y(n_3596)
);

OAI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3423),
.A2(n_1822),
.B(n_1820),
.Y(n_3597)
);

AO21x2_ASAP7_75t_L g3598 ( 
.A1(n_3447),
.A2(n_1828),
.B(n_1824),
.Y(n_3598)
);

AOI21x1_ASAP7_75t_L g3599 ( 
.A1(n_3477),
.A2(n_1833),
.B(n_1829),
.Y(n_3599)
);

INVx5_ASAP7_75t_L g3600 ( 
.A(n_3442),
.Y(n_3600)
);

OAI21x1_ASAP7_75t_L g3601 ( 
.A1(n_3444),
.A2(n_1838),
.B(n_1837),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3479),
.B(n_1853),
.Y(n_3602)
);

OAI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3471),
.A2(n_1841),
.B(n_1840),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3442),
.A2(n_2054),
.B(n_2038),
.Y(n_3604)
);

INVx4_ASAP7_75t_L g3605 ( 
.A(n_3410),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3494),
.A2(n_2054),
.B(n_2439),
.Y(n_3606)
);

A2O1A1Ixp33_ASAP7_75t_L g3607 ( 
.A1(n_3494),
.A2(n_1846),
.B(n_1850),
.C(n_1843),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3458),
.B(n_1555),
.Y(n_3608)
);

BUFx3_ASAP7_75t_L g3609 ( 
.A(n_3507),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3487),
.A2(n_2054),
.B(n_2055),
.Y(n_3610)
);

AOI21x1_ASAP7_75t_SL g3611 ( 
.A1(n_3407),
.A2(n_1558),
.B(n_1556),
.Y(n_3611)
);

AO31x2_ASAP7_75t_L g3612 ( 
.A1(n_3487),
.A2(n_2059),
.A3(n_1860),
.B(n_1867),
.Y(n_3612)
);

INVx3_ASAP7_75t_SL g3613 ( 
.A(n_3466),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3487),
.A2(n_1877),
.B(n_1851),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3424),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3413),
.B(n_1560),
.Y(n_3616)
);

OAI21x1_ASAP7_75t_L g3617 ( 
.A1(n_3487),
.A2(n_1886),
.B(n_1883),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_3417),
.Y(n_3618)
);

OAI22xp5_ASAP7_75t_SL g3619 ( 
.A1(n_3413),
.A2(n_1567),
.B1(n_1572),
.B2(n_1562),
.Y(n_3619)
);

BUFx3_ASAP7_75t_L g3620 ( 
.A(n_3417),
.Y(n_3620)
);

AOI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3413),
.A2(n_1903),
.B(n_1900),
.Y(n_3621)
);

AO21x2_ASAP7_75t_L g3622 ( 
.A1(n_3514),
.A2(n_1912),
.B(n_1910),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3531),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3548),
.Y(n_3624)
);

INVx1_ASAP7_75t_SL g3625 ( 
.A(n_3588),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3544),
.Y(n_3626)
);

AND2x4_ASAP7_75t_L g3627 ( 
.A(n_3574),
.B(n_1013),
.Y(n_3627)
);

OR2x6_ASAP7_75t_L g3628 ( 
.A(n_3582),
.B(n_2838),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3529),
.B(n_1573),
.Y(n_3629)
);

BUFx8_ASAP7_75t_L g3630 ( 
.A(n_3517),
.Y(n_3630)
);

BUFx2_ASAP7_75t_SL g3631 ( 
.A(n_3600),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3561),
.Y(n_3632)
);

BUFx12f_ASAP7_75t_L g3633 ( 
.A(n_3553),
.Y(n_3633)
);

INVx3_ASAP7_75t_SL g3634 ( 
.A(n_3555),
.Y(n_3634)
);

INVx3_ASAP7_75t_L g3635 ( 
.A(n_3523),
.Y(n_3635)
);

OAI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3528),
.A2(n_1576),
.B1(n_1577),
.B2(n_1575),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3510),
.B(n_1579),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_3515),
.B(n_1014),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3615),
.Y(n_3639)
);

AND2x6_ASAP7_75t_L g3640 ( 
.A(n_3620),
.B(n_1919),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3610),
.A2(n_1939),
.B(n_1938),
.Y(n_3641)
);

BUFx2_ASAP7_75t_L g3642 ( 
.A(n_3532),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_3562),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3573),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3512),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3612),
.Y(n_3646)
);

OR2x6_ASAP7_75t_L g3647 ( 
.A(n_3519),
.B(n_2862),
.Y(n_3647)
);

BUFx6f_ASAP7_75t_L g3648 ( 
.A(n_3562),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3550),
.B(n_1016),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3513),
.A2(n_1947),
.B(n_1943),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3554),
.B(n_1580),
.Y(n_3651)
);

INVx5_ASAP7_75t_L g3652 ( 
.A(n_3519),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3525),
.B(n_3621),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3516),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3587),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3590),
.B(n_3575),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3575),
.B(n_1948),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3616),
.B(n_1581),
.Y(n_3658)
);

BUFx12f_ASAP7_75t_L g3659 ( 
.A(n_3605),
.Y(n_3659)
);

INVx2_ASAP7_75t_SL g3660 ( 
.A(n_3537),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3596),
.Y(n_3661)
);

AND2x4_ASAP7_75t_L g3662 ( 
.A(n_3594),
.B(n_1018),
.Y(n_3662)
);

BUFx12f_ASAP7_75t_L g3663 ( 
.A(n_3600),
.Y(n_3663)
);

INVx2_ASAP7_75t_SL g3664 ( 
.A(n_3580),
.Y(n_3664)
);

INVx3_ASAP7_75t_L g3665 ( 
.A(n_3524),
.Y(n_3665)
);

AOI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_3518),
.A2(n_1589),
.B1(n_1590),
.B2(n_1583),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3522),
.A2(n_1958),
.B(n_1957),
.Y(n_3667)
);

INVx5_ASAP7_75t_L g3668 ( 
.A(n_3552),
.Y(n_3668)
);

BUFx3_ASAP7_75t_L g3669 ( 
.A(n_3609),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3577),
.B(n_1591),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3618),
.B(n_1021),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3546),
.B(n_1592),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3549),
.B(n_1594),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_3613),
.Y(n_3674)
);

AND2x4_ASAP7_75t_L g3675 ( 
.A(n_3595),
.B(n_1022),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3612),
.Y(n_3676)
);

HAxp5_ASAP7_75t_L g3677 ( 
.A(n_3560),
.B(n_1853),
.CON(n_3677),
.SN(n_3677)
);

A2O1A1Ixp33_ASAP7_75t_L g3678 ( 
.A1(n_3520),
.A2(n_1964),
.B(n_1965),
.C(n_1959),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3614),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3547),
.B(n_1971),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3572),
.Y(n_3681)
);

BUFx3_ASAP7_75t_L g3682 ( 
.A(n_3591),
.Y(n_3682)
);

HB1xp67_ASAP7_75t_L g3683 ( 
.A(n_3530),
.Y(n_3683)
);

AOI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_3558),
.A2(n_3545),
.B1(n_3597),
.B2(n_3598),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3593),
.B(n_1979),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3538),
.Y(n_3686)
);

INVx3_ASAP7_75t_L g3687 ( 
.A(n_3599),
.Y(n_3687)
);

AND2x4_ASAP7_75t_L g3688 ( 
.A(n_3578),
.B(n_1023),
.Y(n_3688)
);

INVx4_ASAP7_75t_L g3689 ( 
.A(n_3579),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3569),
.A2(n_1604),
.B1(n_1605),
.B2(n_1600),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_L g3691 ( 
.A(n_3535),
.B(n_3559),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3542),
.B(n_1981),
.Y(n_3692)
);

INVx3_ASAP7_75t_L g3693 ( 
.A(n_3564),
.Y(n_3693)
);

INVx5_ASAP7_75t_L g3694 ( 
.A(n_3611),
.Y(n_3694)
);

INVx2_ASAP7_75t_SL g3695 ( 
.A(n_3592),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_3521),
.A2(n_1997),
.B(n_1983),
.Y(n_3696)
);

BUFx6f_ASAP7_75t_L g3697 ( 
.A(n_3608),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3619),
.A2(n_2035),
.B1(n_2041),
.B2(n_1885),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3557),
.Y(n_3699)
);

INVxp67_ASAP7_75t_SL g3700 ( 
.A(n_3576),
.Y(n_3700)
);

BUFx6f_ASAP7_75t_L g3701 ( 
.A(n_3585),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3565),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3567),
.B(n_1999),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3617),
.Y(n_3704)
);

AND2x4_ASAP7_75t_L g3705 ( 
.A(n_3583),
.B(n_1025),
.Y(n_3705)
);

AOI22xp33_ASAP7_75t_L g3706 ( 
.A1(n_3551),
.A2(n_2035),
.B1(n_2041),
.B2(n_1885),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3606),
.B(n_1028),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3581),
.B(n_1607),
.Y(n_3708)
);

HB1xp67_ASAP7_75t_L g3709 ( 
.A(n_3526),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3586),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3511),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3540),
.Y(n_3712)
);

AND2x4_ASAP7_75t_L g3713 ( 
.A(n_3601),
.B(n_1036),
.Y(n_3713)
);

INVx5_ASAP7_75t_L g3714 ( 
.A(n_3607),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3511),
.Y(n_3715)
);

NAND2x1_ASAP7_75t_L g3716 ( 
.A(n_3536),
.B(n_2001),
.Y(n_3716)
);

AND2x4_ASAP7_75t_L g3717 ( 
.A(n_3642),
.B(n_3584),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3645),
.B(n_3603),
.Y(n_3718)
);

OAI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3696),
.A2(n_3715),
.B(n_3676),
.Y(n_3719)
);

OAI21x1_ASAP7_75t_L g3720 ( 
.A1(n_3646),
.A2(n_3533),
.B(n_3571),
.Y(n_3720)
);

NAND3xp33_ASAP7_75t_L g3721 ( 
.A(n_3666),
.B(n_3589),
.C(n_3534),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3700),
.B(n_3570),
.Y(n_3722)
);

BUFx3_ASAP7_75t_L g3723 ( 
.A(n_3652),
.Y(n_3723)
);

CKINVDCx5p33_ASAP7_75t_R g3724 ( 
.A(n_3633),
.Y(n_3724)
);

AND2x4_ASAP7_75t_L g3725 ( 
.A(n_3682),
.B(n_3604),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3626),
.Y(n_3726)
);

OA21x2_ASAP7_75t_L g3727 ( 
.A1(n_3667),
.A2(n_3541),
.B(n_3563),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3632),
.Y(n_3728)
);

BUFx6f_ASAP7_75t_L g3729 ( 
.A(n_3663),
.Y(n_3729)
);

OAI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3653),
.A2(n_3539),
.B(n_3566),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3639),
.Y(n_3731)
);

NOR2xp67_ASAP7_75t_L g3732 ( 
.A(n_3668),
.B(n_3543),
.Y(n_3732)
);

OR3x4_ASAP7_75t_SL g3733 ( 
.A(n_3630),
.B(n_3634),
.C(n_3677),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3711),
.A2(n_3527),
.B(n_3556),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3704),
.A2(n_3568),
.B(n_2005),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3625),
.B(n_3602),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3684),
.A2(n_1613),
.B1(n_1614),
.B2(n_1608),
.Y(n_3737)
);

AOI22x1_ASAP7_75t_L g3738 ( 
.A1(n_3650),
.A2(n_1616),
.B1(n_1617),
.B2(n_1615),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3644),
.B(n_1622),
.Y(n_3739)
);

OAI21x1_ASAP7_75t_SL g3740 ( 
.A1(n_3712),
.A2(n_2010),
.B(n_2003),
.Y(n_3740)
);

AO21x2_ASAP7_75t_L g3741 ( 
.A1(n_3686),
.A2(n_2014),
.B(n_2013),
.Y(n_3741)
);

BUFx5_ASAP7_75t_L g3742 ( 
.A(n_3702),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3661),
.Y(n_3743)
);

INVx2_ASAP7_75t_SL g3744 ( 
.A(n_3652),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3693),
.A2(n_2034),
.B(n_2027),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3699),
.A2(n_2044),
.B(n_2761),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3655),
.Y(n_3747)
);

INVxp67_ASAP7_75t_L g3748 ( 
.A(n_3695),
.Y(n_3748)
);

OAI21x1_ASAP7_75t_L g3749 ( 
.A1(n_3710),
.A2(n_2836),
.B(n_1038),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3643),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3654),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3624),
.Y(n_3752)
);

OAI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3714),
.A2(n_1624),
.B1(n_1625),
.B2(n_1623),
.Y(n_3753)
);

AOI221xp5_ASAP7_75t_L g3754 ( 
.A1(n_3685),
.A2(n_1633),
.B1(n_1635),
.B2(n_1631),
.C(n_1626),
.Y(n_3754)
);

OAI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3681),
.A2(n_1041),
.B(n_1037),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3691),
.A2(n_1641),
.B1(n_1642),
.B2(n_1638),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3679),
.A2(n_1045),
.B(n_1044),
.Y(n_3757)
);

AOI22xp33_ASAP7_75t_L g3758 ( 
.A1(n_3714),
.A2(n_1645),
.B1(n_1647),
.B2(n_1644),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_L g3759 ( 
.A(n_3651),
.B(n_1648),
.Y(n_3759)
);

OAI21x1_ASAP7_75t_L g3760 ( 
.A1(n_3687),
.A2(n_1051),
.B(n_1048),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_SL g3761 ( 
.A(n_3659),
.B(n_1651),
.Y(n_3761)
);

OAI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3683),
.A2(n_1054),
.B(n_1052),
.Y(n_3762)
);

OAI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3706),
.A2(n_1658),
.B(n_1656),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3656),
.A2(n_1665),
.B(n_1663),
.Y(n_3764)
);

OA21x2_ASAP7_75t_L g3765 ( 
.A1(n_3678),
.A2(n_1674),
.B(n_1666),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3709),
.A2(n_3622),
.B(n_3628),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3623),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_SL g3768 ( 
.A1(n_3637),
.A2(n_1683),
.B(n_1677),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3657),
.Y(n_3769)
);

OAI21x1_ASAP7_75t_L g3770 ( 
.A1(n_3641),
.A2(n_1056),
.B(n_1055),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_SL g3771 ( 
.A(n_3694),
.B(n_1684),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3716),
.A2(n_3680),
.B(n_3692),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3665),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_3648),
.Y(n_3774)
);

BUFx2_ASAP7_75t_L g3775 ( 
.A(n_3674),
.Y(n_3775)
);

INVxp67_ASAP7_75t_L g3776 ( 
.A(n_3664),
.Y(n_3776)
);

BUFx6f_ASAP7_75t_L g3777 ( 
.A(n_3669),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3694),
.A2(n_1687),
.B(n_1685),
.Y(n_3778)
);

OA21x2_ASAP7_75t_L g3779 ( 
.A1(n_3705),
.A2(n_1692),
.B(n_1691),
.Y(n_3779)
);

OR2x2_ASAP7_75t_L g3780 ( 
.A(n_3670),
.B(n_2),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3689),
.Y(n_3781)
);

AND2x4_ASAP7_75t_L g3782 ( 
.A(n_3635),
.B(n_1057),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_L g3783 ( 
.A1(n_3703),
.A2(n_1059),
.B(n_1058),
.Y(n_3783)
);

OA21x2_ASAP7_75t_L g3784 ( 
.A1(n_3713),
.A2(n_1698),
.B(n_1696),
.Y(n_3784)
);

OAI21x1_ASAP7_75t_L g3785 ( 
.A1(n_3629),
.A2(n_1063),
.B(n_1060),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3631),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3658),
.A2(n_3673),
.B(n_3672),
.Y(n_3787)
);

INVx2_ASAP7_75t_SL g3788 ( 
.A(n_3660),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3640),
.A2(n_3701),
.B1(n_3707),
.B2(n_3697),
.Y(n_3789)
);

AO31x2_ASAP7_75t_L g3790 ( 
.A1(n_3636),
.A2(n_4),
.A3(n_2),
.B(n_3),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3675),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3638),
.Y(n_3792)
);

INVx4_ASAP7_75t_L g3793 ( 
.A(n_3777),
.Y(n_3793)
);

AND2x4_ASAP7_75t_L g3794 ( 
.A(n_3775),
.B(n_3627),
.Y(n_3794)
);

OR2x6_ASAP7_75t_L g3795 ( 
.A(n_3766),
.B(n_3671),
.Y(n_3795)
);

INVx3_ASAP7_75t_L g3796 ( 
.A(n_3777),
.Y(n_3796)
);

AND2x4_ASAP7_75t_L g3797 ( 
.A(n_3751),
.B(n_3662),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3750),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_L g3799 ( 
.A1(n_3721),
.A2(n_3640),
.B1(n_3688),
.B2(n_3698),
.Y(n_3799)
);

AND2x2_ASAP7_75t_SL g3800 ( 
.A(n_3784),
.B(n_3649),
.Y(n_3800)
);

INVx1_ASAP7_75t_SL g3801 ( 
.A(n_3736),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3747),
.B(n_3708),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3720),
.A2(n_3690),
.B(n_1067),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3743),
.B(n_1699),
.Y(n_3804)
);

AND2x2_ASAP7_75t_SL g3805 ( 
.A(n_3779),
.B(n_3647),
.Y(n_3805)
);

AOI222xp33_ASAP7_75t_L g3806 ( 
.A1(n_3754),
.A2(n_1705),
.B1(n_1701),
.B2(n_1707),
.C1(n_1703),
.C2(n_1700),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_3774),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3764),
.A2(n_1715),
.B1(n_1717),
.B2(n_1708),
.Y(n_3808)
);

BUFx10_ASAP7_75t_L g3809 ( 
.A(n_3724),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3759),
.A2(n_1722),
.B1(n_1727),
.B2(n_1719),
.Y(n_3810)
);

INVx3_ASAP7_75t_L g3811 ( 
.A(n_3723),
.Y(n_3811)
);

HB1xp67_ASAP7_75t_L g3812 ( 
.A(n_3781),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3728),
.B(n_1066),
.Y(n_3813)
);

AO21x2_ASAP7_75t_L g3814 ( 
.A1(n_3740),
.A2(n_3),
.B(n_4),
.Y(n_3814)
);

NAND2x1p5_ASAP7_75t_L g3815 ( 
.A(n_3717),
.B(n_2862),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_SL g3816 ( 
.A1(n_3765),
.A2(n_3730),
.B1(n_3741),
.B2(n_3722),
.Y(n_3816)
);

BUFx3_ASAP7_75t_L g3817 ( 
.A(n_3729),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3737),
.A2(n_2039),
.B(n_2042),
.C(n_2036),
.Y(n_3818)
);

BUFx12f_ASAP7_75t_L g3819 ( 
.A(n_3729),
.Y(n_3819)
);

NAND2xp33_ASAP7_75t_L g3820 ( 
.A(n_3758),
.B(n_1729),
.Y(n_3820)
);

AND2x2_ASAP7_75t_SL g3821 ( 
.A(n_3769),
.B(n_6),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3726),
.B(n_3731),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3738),
.A2(n_1732),
.B1(n_1733),
.B2(n_1730),
.Y(n_3823)
);

HB1xp67_ASAP7_75t_L g3824 ( 
.A(n_3767),
.Y(n_3824)
);

AOI22xp33_ASAP7_75t_L g3825 ( 
.A1(n_3725),
.A2(n_1736),
.B1(n_1740),
.B2(n_1734),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3748),
.B(n_1741),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3792),
.A2(n_1745),
.B1(n_1746),
.B2(n_1744),
.Y(n_3827)
);

INVx2_ASAP7_75t_SL g3828 ( 
.A(n_3788),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3752),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_3789),
.B(n_1748),
.Y(n_3830)
);

CKINVDCx14_ASAP7_75t_R g3831 ( 
.A(n_3780),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_SL g3832 ( 
.A1(n_3744),
.A2(n_1752),
.B1(n_1755),
.B2(n_1751),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3791),
.A2(n_1759),
.B1(n_1767),
.B2(n_1757),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3742),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3742),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3786),
.B(n_7),
.Y(n_3836)
);

AOI22xp33_ASAP7_75t_SL g3837 ( 
.A1(n_3753),
.A2(n_3772),
.B1(n_3787),
.B2(n_3783),
.Y(n_3837)
);

INVx2_ASAP7_75t_SL g3838 ( 
.A(n_3773),
.Y(n_3838)
);

INVx4_ASAP7_75t_L g3839 ( 
.A(n_3733),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_SL g3840 ( 
.A1(n_3785),
.A2(n_1772),
.B1(n_1773),
.B2(n_1770),
.Y(n_3840)
);

OAI22xp33_ASAP7_75t_L g3841 ( 
.A1(n_3718),
.A2(n_1775),
.B1(n_1777),
.B2(n_1774),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3734),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3742),
.Y(n_3843)
);

INVx3_ASAP7_75t_L g3844 ( 
.A(n_3782),
.Y(n_3844)
);

AOI221xp5_ASAP7_75t_L g3845 ( 
.A1(n_3756),
.A2(n_2016),
.B1(n_2018),
.B2(n_2015),
.C(n_2011),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3719),
.Y(n_3846)
);

OAI221xp5_ASAP7_75t_L g3847 ( 
.A1(n_3768),
.A2(n_1791),
.B1(n_1794),
.B2(n_1779),
.C(n_1778),
.Y(n_3847)
);

OAI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3732),
.A2(n_2053),
.B1(n_2058),
.B2(n_2049),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3790),
.Y(n_3849)
);

NOR2xp67_ASAP7_75t_L g3850 ( 
.A(n_3776),
.B(n_8),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3790),
.Y(n_3851)
);

OR2x2_ASAP7_75t_L g3852 ( 
.A(n_3739),
.B(n_9),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3735),
.B(n_1796),
.Y(n_3853)
);

NAND2x1_ASAP7_75t_L g3854 ( 
.A(n_3727),
.B(n_9),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3771),
.B(n_3745),
.Y(n_3855)
);

AOI22xp33_ASAP7_75t_SL g3856 ( 
.A1(n_3762),
.A2(n_1802),
.B1(n_1805),
.B2(n_1799),
.Y(n_3856)
);

INVx3_ASAP7_75t_L g3857 ( 
.A(n_3755),
.Y(n_3857)
);

INVx1_ASAP7_75t_SL g3858 ( 
.A(n_3761),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3746),
.B(n_10),
.Y(n_3859)
);

OAI21x1_ASAP7_75t_L g3860 ( 
.A1(n_3749),
.A2(n_1073),
.B(n_1072),
.Y(n_3860)
);

AOI22xp5_ASAP7_75t_L g3861 ( 
.A1(n_3770),
.A2(n_1809),
.B1(n_1811),
.B2(n_1806),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3757),
.Y(n_3862)
);

AOI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_3763),
.A2(n_1825),
.B1(n_1826),
.B2(n_1812),
.Y(n_3863)
);

NAND2x1p5_ASAP7_75t_L g3864 ( 
.A(n_3760),
.B(n_3778),
.Y(n_3864)
);

INVx2_ASAP7_75t_SL g3865 ( 
.A(n_3777),
.Y(n_3865)
);

CKINVDCx20_ASAP7_75t_R g3866 ( 
.A(n_3724),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3726),
.Y(n_3867)
);

BUFx6f_ASAP7_75t_L g3868 ( 
.A(n_3777),
.Y(n_3868)
);

AOI22xp5_ASAP7_75t_L g3869 ( 
.A1(n_3721),
.A2(n_1832),
.B1(n_1836),
.B2(n_1827),
.Y(n_3869)
);

OAI21x1_ASAP7_75t_L g3870 ( 
.A1(n_3854),
.A2(n_10),
.B(n_11),
.Y(n_3870)
);

AOI21x1_ASAP7_75t_L g3871 ( 
.A1(n_3855),
.A2(n_1842),
.B(n_1839),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3867),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3812),
.Y(n_3873)
);

OA21x2_ASAP7_75t_L g3874 ( 
.A1(n_3834),
.A2(n_1852),
.B(n_1844),
.Y(n_3874)
);

INVx2_ASAP7_75t_SL g3875 ( 
.A(n_3868),
.Y(n_3875)
);

BUFx3_ASAP7_75t_L g3876 ( 
.A(n_3819),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3838),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3824),
.Y(n_3878)
);

AND2x4_ASAP7_75t_L g3879 ( 
.A(n_3811),
.B(n_11),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3822),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3829),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3849),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3835),
.Y(n_3883)
);

AOI21x1_ASAP7_75t_L g3884 ( 
.A1(n_3851),
.A2(n_1856),
.B(n_1854),
.Y(n_3884)
);

INVx5_ASAP7_75t_L g3885 ( 
.A(n_3839),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3801),
.B(n_12),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3843),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3842),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3846),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_3793),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3802),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3862),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3828),
.Y(n_3893)
);

OR2x2_ASAP7_75t_L g3894 ( 
.A(n_3804),
.B(n_13),
.Y(n_3894)
);

INVx4_ASAP7_75t_L g3895 ( 
.A(n_3868),
.Y(n_3895)
);

BUFx3_ASAP7_75t_L g3896 ( 
.A(n_3866),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3857),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3836),
.Y(n_3898)
);

INVx2_ASAP7_75t_SL g3899 ( 
.A(n_3796),
.Y(n_3899)
);

INVx1_ASAP7_75t_SL g3900 ( 
.A(n_3807),
.Y(n_3900)
);

INVx2_ASAP7_75t_SL g3901 ( 
.A(n_3865),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3798),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3797),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3795),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3816),
.A2(n_1866),
.B(n_1859),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3831),
.B(n_1868),
.Y(n_3906)
);

AND2x4_ASAP7_75t_L g3907 ( 
.A(n_3794),
.B(n_13),
.Y(n_3907)
);

BUFx3_ASAP7_75t_L g3908 ( 
.A(n_3817),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3859),
.Y(n_3909)
);

CKINVDCx5p33_ASAP7_75t_R g3910 ( 
.A(n_3809),
.Y(n_3910)
);

AO21x2_ASAP7_75t_L g3911 ( 
.A1(n_3853),
.A2(n_14),
.B(n_15),
.Y(n_3911)
);

OAI21x1_ASAP7_75t_L g3912 ( 
.A1(n_3803),
.A2(n_17),
.B(n_18),
.Y(n_3912)
);

INVx3_ASAP7_75t_L g3913 ( 
.A(n_3798),
.Y(n_3913)
);

INVx2_ASAP7_75t_SL g3914 ( 
.A(n_3844),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3795),
.B(n_18),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3815),
.Y(n_3916)
);

BUFx2_ASAP7_75t_L g3917 ( 
.A(n_3800),
.Y(n_3917)
);

INVx2_ASAP7_75t_SL g3918 ( 
.A(n_3826),
.Y(n_3918)
);

AO21x2_ASAP7_75t_L g3919 ( 
.A1(n_3850),
.A2(n_19),
.B(n_21),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3858),
.B(n_19),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3852),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3814),
.Y(n_3922)
);

INVx4_ASAP7_75t_L g3923 ( 
.A(n_3813),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3837),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3805),
.B(n_21),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3821),
.Y(n_3926)
);

AOI22xp33_ASAP7_75t_L g3927 ( 
.A1(n_3799),
.A2(n_1990),
.B1(n_1991),
.B2(n_1988),
.Y(n_3927)
);

HB1xp67_ASAP7_75t_L g3928 ( 
.A(n_3864),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3860),
.Y(n_3929)
);

INVx3_ASAP7_75t_L g3930 ( 
.A(n_3830),
.Y(n_3930)
);

OAI21x1_ASAP7_75t_L g3931 ( 
.A1(n_3861),
.A2(n_22),
.B(n_23),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3833),
.B(n_22),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3869),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3827),
.Y(n_3934)
);

INVx3_ASAP7_75t_L g3935 ( 
.A(n_3848),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3832),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3882),
.Y(n_3937)
);

AOI221xp5_ASAP7_75t_L g3938 ( 
.A1(n_3905),
.A2(n_3841),
.B1(n_3847),
.B2(n_3810),
.C(n_3808),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3872),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_SL g3940 ( 
.A1(n_3924),
.A2(n_3820),
.B1(n_3840),
.B2(n_3856),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3881),
.Y(n_3941)
);

AOI221xp5_ASAP7_75t_L g3942 ( 
.A1(n_3933),
.A2(n_3845),
.B1(n_3818),
.B2(n_1873),
.C(n_1875),
.Y(n_3942)
);

OAI211xp5_ASAP7_75t_L g3943 ( 
.A1(n_3927),
.A2(n_3863),
.B(n_3806),
.C(n_3825),
.Y(n_3943)
);

OAI211xp5_ASAP7_75t_SL g3944 ( 
.A1(n_3935),
.A2(n_3934),
.B(n_3909),
.C(n_3921),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_SL g3945 ( 
.A(n_3876),
.Y(n_3945)
);

INVxp67_ASAP7_75t_L g3946 ( 
.A(n_3891),
.Y(n_3946)
);

AO21x2_ASAP7_75t_L g3947 ( 
.A1(n_3922),
.A2(n_23),
.B(n_24),
.Y(n_3947)
);

OAI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3917),
.A2(n_3823),
.B1(n_1871),
.B2(n_1878),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_SL g3949 ( 
.A1(n_3930),
.A2(n_3925),
.B1(n_3911),
.B2(n_3874),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3936),
.A2(n_1880),
.B1(n_1887),
.B2(n_1870),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3889),
.Y(n_3951)
);

AOI22xp33_ASAP7_75t_L g3952 ( 
.A1(n_3904),
.A2(n_1890),
.B1(n_1891),
.B2(n_1888),
.Y(n_3952)
);

OAI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3926),
.A2(n_1894),
.B1(n_1895),
.B2(n_1892),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3883),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3885),
.A2(n_1898),
.B1(n_1899),
.B2(n_1897),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3914),
.B(n_3903),
.Y(n_3956)
);

AND2x4_ASAP7_75t_L g3957 ( 
.A(n_3916),
.B(n_3877),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3918),
.A2(n_1905),
.B1(n_1909),
.B2(n_1904),
.Y(n_3958)
);

OAI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3900),
.A2(n_3899),
.B1(n_3885),
.B2(n_3893),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3929),
.A2(n_1916),
.B1(n_1922),
.B2(n_1915),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3888),
.Y(n_3961)
);

OAI21xp5_ASAP7_75t_SL g3962 ( 
.A1(n_3871),
.A2(n_34),
.B(n_25),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_L g3963 ( 
.A1(n_3931),
.A2(n_3932),
.B1(n_3928),
.B2(n_3923),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3880),
.Y(n_3964)
);

OAI21x1_ASAP7_75t_L g3965 ( 
.A1(n_3897),
.A2(n_25),
.B(n_27),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3915),
.A2(n_1925),
.B1(n_1926),
.B2(n_1924),
.Y(n_3966)
);

OAI22xp33_ASAP7_75t_L g3967 ( 
.A1(n_3886),
.A2(n_1930),
.B1(n_1932),
.B2(n_1927),
.Y(n_3967)
);

OAI211xp5_ASAP7_75t_L g3968 ( 
.A1(n_3884),
.A2(n_1937),
.B(n_1940),
.C(n_1935),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3898),
.A2(n_1949),
.B1(n_1951),
.B2(n_1946),
.Y(n_3969)
);

A2O1A1Ixp33_ASAP7_75t_L g3970 ( 
.A1(n_3870),
.A2(n_1984),
.B(n_2047),
.C(n_1968),
.Y(n_3970)
);

OR2x2_ASAP7_75t_L g3971 ( 
.A(n_3878),
.B(n_28),
.Y(n_3971)
);

AND2x2_ASAP7_75t_SL g3972 ( 
.A(n_3879),
.B(n_29),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3887),
.Y(n_3973)
);

AOI21x1_ASAP7_75t_L g3974 ( 
.A1(n_3906),
.A2(n_1960),
.B(n_1955),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3919),
.A2(n_1969),
.B1(n_1970),
.B2(n_1967),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3894),
.A2(n_1973),
.B1(n_1974),
.B2(n_1972),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3873),
.B(n_29),
.Y(n_3977)
);

AOI22xp33_ASAP7_75t_L g3978 ( 
.A1(n_3890),
.A2(n_1977),
.B1(n_1992),
.B2(n_1976),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3892),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3901),
.Y(n_3980)
);

OAI211xp5_ASAP7_75t_SL g3981 ( 
.A1(n_3902),
.A2(n_1995),
.B(n_2004),
.C(n_1993),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3913),
.B(n_3875),
.Y(n_3982)
);

AND2x4_ASAP7_75t_L g3983 ( 
.A(n_3908),
.B(n_30),
.Y(n_3983)
);

OAI22xp5_ASAP7_75t_L g3984 ( 
.A1(n_3895),
.A2(n_3907),
.B1(n_3910),
.B2(n_3896),
.Y(n_3984)
);

AOI22xp5_ASAP7_75t_L g3985 ( 
.A1(n_3920),
.A2(n_2026),
.B1(n_2030),
.B2(n_2008),
.Y(n_3985)
);

AOI22xp33_ASAP7_75t_L g3986 ( 
.A1(n_3912),
.A2(n_2060),
.B1(n_2061),
.B2(n_2048),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3883),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3888),
.Y(n_3988)
);

OAI211xp5_ASAP7_75t_L g3989 ( 
.A1(n_3905),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_3989)
);

BUFx6f_ASAP7_75t_L g3990 ( 
.A(n_3876),
.Y(n_3990)
);

AOI22xp33_ASAP7_75t_L g3991 ( 
.A1(n_3924),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3883),
.Y(n_3992)
);

AOI21x1_ASAP7_75t_L g3993 ( 
.A1(n_3925),
.A2(n_35),
.B(n_36),
.Y(n_3993)
);

HB1xp67_ASAP7_75t_L g3994 ( 
.A(n_3888),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_SL g3995 ( 
.A1(n_3924),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_3995)
);

OA21x2_ASAP7_75t_L g3996 ( 
.A1(n_3924),
.A2(n_38),
.B(n_39),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3895),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3883),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3882),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3891),
.B(n_38),
.Y(n_4000)
);

OA21x2_ASAP7_75t_L g4001 ( 
.A1(n_3924),
.A2(n_40),
.B(n_41),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3882),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3891),
.B(n_41),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3883),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_SL g4005 ( 
.A(n_3924),
.B(n_43),
.C(n_44),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3882),
.Y(n_4006)
);

OAI221xp5_ASAP7_75t_L g4007 ( 
.A1(n_3905),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3909),
.B(n_46),
.Y(n_4008)
);

INVx2_ASAP7_75t_SL g4009 ( 
.A(n_3908),
.Y(n_4009)
);

OAI332xp33_ASAP7_75t_L g4010 ( 
.A1(n_3933),
.A2(n_52),
.A3(n_51),
.B1(n_49),
.B2(n_53),
.B3(n_47),
.C1(n_48),
.C2(n_50),
.Y(n_4010)
);

OAI21xp33_ASAP7_75t_L g4011 ( 
.A1(n_3924),
.A2(n_51),
.B(n_50),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3882),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3882),
.Y(n_4013)
);

INVx11_ASAP7_75t_L g4014 ( 
.A(n_3896),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3924),
.A2(n_54),
.B1(n_48),
.B2(n_53),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3883),
.Y(n_4016)
);

A2O1A1Ixp33_ASAP7_75t_L g4017 ( 
.A1(n_3905),
.A2(n_63),
.B(n_71),
.C(n_54),
.Y(n_4017)
);

NAND3xp33_ASAP7_75t_L g4018 ( 
.A(n_3905),
.B(n_55),
.C(n_56),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3891),
.B(n_55),
.Y(n_4019)
);

AOI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3924),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3882),
.Y(n_4021)
);

HB1xp67_ASAP7_75t_L g4022 ( 
.A(n_3888),
.Y(n_4022)
);

OAI221xp5_ASAP7_75t_SL g4023 ( 
.A1(n_3927),
.A2(n_60),
.B1(n_57),
.B2(n_58),
.C(n_61),
.Y(n_4023)
);

OAI21x1_ASAP7_75t_L g4024 ( 
.A1(n_3882),
.A2(n_60),
.B(n_61),
.Y(n_4024)
);

AND2x4_ASAP7_75t_SL g4025 ( 
.A(n_3895),
.B(n_63),
.Y(n_4025)
);

OAI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3924),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_4026)
);

OA21x2_ASAP7_75t_L g4027 ( 
.A1(n_3924),
.A2(n_64),
.B(n_65),
.Y(n_4027)
);

OR2x2_ASAP7_75t_L g4028 ( 
.A(n_3909),
.B(n_67),
.Y(n_4028)
);

AOI221xp5_ASAP7_75t_L g4029 ( 
.A1(n_3905),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_4029)
);

AOI222xp33_ASAP7_75t_L g4030 ( 
.A1(n_3905),
.A2(n_70),
.B1(n_73),
.B2(n_68),
.C1(n_69),
.C2(n_72),
.Y(n_4030)
);

OAI221xp5_ASAP7_75t_L g4031 ( 
.A1(n_3905),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.C(n_76),
.Y(n_4031)
);

OAI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3924),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_4032)
);

INVx3_ASAP7_75t_L g4033 ( 
.A(n_3895),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3924),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_4034)
);

OR2x2_ASAP7_75t_L g4035 ( 
.A(n_3909),
.B(n_77),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3917),
.B(n_80),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3882),
.Y(n_4037)
);

AOI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3924),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3882),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3924),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_4040)
);

OAI22xp33_ASAP7_75t_L g4041 ( 
.A1(n_3924),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4041)
);

OA21x2_ASAP7_75t_L g4042 ( 
.A1(n_3924),
.A2(n_86),
.B(n_87),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3924),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3924),
.A2(n_88),
.B(n_89),
.Y(n_4044)
);

INVx5_ASAP7_75t_SL g4045 ( 
.A(n_3919),
.Y(n_4045)
);

OA21x2_ASAP7_75t_L g4046 ( 
.A1(n_3924),
.A2(n_90),
.B(n_91),
.Y(n_4046)
);

OAI221xp5_ASAP7_75t_L g4047 ( 
.A1(n_3905),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.C(n_95),
.Y(n_4047)
);

O2A1O1Ixp33_ASAP7_75t_SL g4048 ( 
.A1(n_3926),
.A2(n_95),
.B(n_92),
.C(n_93),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3882),
.Y(n_4049)
);

AO21x2_ASAP7_75t_L g4050 ( 
.A1(n_3922),
.A2(n_96),
.B(n_97),
.Y(n_4050)
);

AO22x2_ASAP7_75t_L g4051 ( 
.A1(n_3924),
.A2(n_98),
.B1(n_99),
.B2(n_97),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3924),
.A2(n_100),
.B1(n_96),
.B2(n_98),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_3924),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3882),
.Y(n_4054)
);

AND2x4_ASAP7_75t_L g4055 ( 
.A(n_3997),
.B(n_101),
.Y(n_4055)
);

OR2x2_ASAP7_75t_L g4056 ( 
.A(n_3946),
.B(n_102),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3982),
.B(n_3956),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3980),
.B(n_4033),
.Y(n_4058)
);

OR2x2_ASAP7_75t_L g4059 ( 
.A(n_3964),
.B(n_103),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3959),
.B(n_104),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3954),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3957),
.B(n_104),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3987),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3992),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3937),
.Y(n_4065)
);

OR2x2_ASAP7_75t_L g4066 ( 
.A(n_3939),
.B(n_105),
.Y(n_4066)
);

BUFx3_ASAP7_75t_L g4067 ( 
.A(n_3990),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_3963),
.B(n_105),
.Y(n_4068)
);

OR2x2_ASAP7_75t_L g4069 ( 
.A(n_3971),
.B(n_106),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_4009),
.B(n_106),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_3998),
.B(n_107),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_3973),
.B(n_108),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_3961),
.B(n_108),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3999),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_4002),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_4004),
.B(n_109),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_4006),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4012),
.Y(n_4078)
);

OR2x2_ASAP7_75t_L g4079 ( 
.A(n_3988),
.B(n_109),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_3994),
.B(n_4022),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_SL g4081 ( 
.A1(n_4045),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_3951),
.Y(n_4082)
);

OR2x2_ASAP7_75t_L g4083 ( 
.A(n_3941),
.B(n_112),
.Y(n_4083)
);

BUFx2_ASAP7_75t_L g4084 ( 
.A(n_3996),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4013),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4021),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_4016),
.Y(n_4087)
);

NOR2xp67_ASAP7_75t_L g4088 ( 
.A(n_3984),
.B(n_114),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4037),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3979),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_4036),
.B(n_3977),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3940),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4092)
);

OR2x2_ASAP7_75t_SL g4093 ( 
.A(n_4001),
.B(n_116),
.Y(n_4093)
);

INVx4_ASAP7_75t_L g4094 ( 
.A(n_3990),
.Y(n_4094)
);

OR2x2_ASAP7_75t_L g4095 ( 
.A(n_4008),
.B(n_115),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_4039),
.B(n_117),
.Y(n_4096)
);

AND2x4_ASAP7_75t_L g4097 ( 
.A(n_4028),
.B(n_4035),
.Y(n_4097)
);

INVx1_ASAP7_75t_SL g4098 ( 
.A(n_4025),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4049),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3949),
.B(n_118),
.Y(n_4100)
);

HB1xp67_ASAP7_75t_L g4101 ( 
.A(n_4054),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_SL g4102 ( 
.A1(n_4045),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4000),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_4003),
.B(n_119),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_4018),
.A2(n_124),
.B1(n_120),
.B2(n_122),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_4027),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_4019),
.B(n_122),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_4042),
.B(n_124),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3947),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4046),
.B(n_125),
.Y(n_4110)
);

INVx2_ASAP7_75t_SL g4111 ( 
.A(n_4014),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4050),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4024),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4051),
.B(n_126),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3965),
.Y(n_4115)
);

AND2x2_ASAP7_75t_L g4116 ( 
.A(n_3972),
.B(n_127),
.Y(n_4116)
);

AND2x4_ASAP7_75t_L g4117 ( 
.A(n_3983),
.B(n_128),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_4051),
.B(n_128),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3993),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3945),
.Y(n_4120)
);

NOR2xp33_ASAP7_75t_L g4121 ( 
.A(n_3974),
.B(n_129),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3967),
.B(n_130),
.Y(n_4122)
);

HB1xp67_ASAP7_75t_L g4123 ( 
.A(n_4015),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_4026),
.Y(n_4124)
);

AOI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_4007),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3944),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4034),
.Y(n_4127)
);

INVx3_ASAP7_75t_L g4128 ( 
.A(n_4005),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_4044),
.B(n_131),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_3985),
.B(n_133),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_3962),
.Y(n_4131)
);

INVx2_ASAP7_75t_SL g4132 ( 
.A(n_3948),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_3955),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_3976),
.B(n_134),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3966),
.B(n_3952),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_4031),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4136)
);

BUFx3_ASAP7_75t_L g4137 ( 
.A(n_4047),
.Y(n_4137)
);

AND3x2_ASAP7_75t_L g4138 ( 
.A(n_4029),
.B(n_135),
.C(n_137),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4011),
.B(n_138),
.Y(n_4139)
);

BUFx2_ASAP7_75t_SL g4140 ( 
.A(n_4048),
.Y(n_4140)
);

CKINVDCx20_ASAP7_75t_R g4141 ( 
.A(n_3943),
.Y(n_4141)
);

AND2x4_ASAP7_75t_L g4142 ( 
.A(n_3970),
.B(n_138),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4032),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_3969),
.B(n_139),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_3986),
.B(n_3995),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4041),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3975),
.B(n_139),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3953),
.B(n_140),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3991),
.B(n_140),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4020),
.B(n_142),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4038),
.B(n_143),
.Y(n_4151)
);

INVx2_ASAP7_75t_SL g4152 ( 
.A(n_4010),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3968),
.Y(n_4153)
);

INVxp67_ASAP7_75t_L g4154 ( 
.A(n_4030),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4040),
.Y(n_4155)
);

INVxp67_ASAP7_75t_SL g4156 ( 
.A(n_4053),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_4043),
.B(n_143),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4052),
.Y(n_4158)
);

HB1xp67_ASAP7_75t_L g4159 ( 
.A(n_3989),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3950),
.B(n_145),
.Y(n_4160)
);

AOI22xp33_ASAP7_75t_L g4161 ( 
.A1(n_3938),
.A2(n_148),
.B1(n_145),
.B2(n_146),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3960),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4017),
.Y(n_4163)
);

OR2x2_ASAP7_75t_L g4164 ( 
.A(n_3958),
.B(n_146),
.Y(n_4164)
);

OR2x2_ASAP7_75t_L g4165 ( 
.A(n_4023),
.B(n_148),
.Y(n_4165)
);

AND2x4_ASAP7_75t_SL g4166 ( 
.A(n_3978),
.B(n_149),
.Y(n_4166)
);

AND2x4_ASAP7_75t_L g4167 ( 
.A(n_3981),
.B(n_150),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3942),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3954),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3946),
.B(n_150),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3937),
.Y(n_4171)
);

BUFx6f_ASAP7_75t_L g4172 ( 
.A(n_3990),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3946),
.B(n_151),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3946),
.B(n_151),
.Y(n_4174)
);

HB1xp67_ASAP7_75t_L g4175 ( 
.A(n_3961),
.Y(n_4175)
);

AND2x4_ASAP7_75t_SL g4176 ( 
.A(n_3990),
.B(n_152),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_3946),
.B(n_152),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3946),
.B(n_153),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_3982),
.B(n_153),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3946),
.B(n_154),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_3982),
.B(n_154),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3937),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3946),
.B(n_155),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3937),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3937),
.Y(n_4185)
);

AND2x4_ASAP7_75t_L g4186 ( 
.A(n_3997),
.B(n_155),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3937),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_SL g4188 ( 
.A(n_3949),
.B(n_156),
.Y(n_4188)
);

BUFx2_ASAP7_75t_L g4189 ( 
.A(n_3997),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3937),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3937),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_3982),
.B(n_157),
.Y(n_4192)
);

BUFx2_ASAP7_75t_L g4193 ( 
.A(n_3997),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3937),
.Y(n_4194)
);

HB1xp67_ASAP7_75t_L g4195 ( 
.A(n_3961),
.Y(n_4195)
);

OR2x2_ASAP7_75t_L g4196 ( 
.A(n_3946),
.B(n_157),
.Y(n_4196)
);

NOR2x1p5_ASAP7_75t_L g4197 ( 
.A(n_4005),
.B(n_158),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3946),
.B(n_158),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3937),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3937),
.Y(n_4200)
);

OR2x2_ASAP7_75t_L g4201 ( 
.A(n_3946),
.B(n_159),
.Y(n_4201)
);

INVx5_ASAP7_75t_L g4202 ( 
.A(n_3990),
.Y(n_4202)
);

INVxp67_ASAP7_75t_SL g4203 ( 
.A(n_3996),
.Y(n_4203)
);

BUFx2_ASAP7_75t_L g4204 ( 
.A(n_3997),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3946),
.B(n_159),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3937),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_3946),
.B(n_161),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3940),
.A2(n_164),
.B1(n_161),
.B2(n_163),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3937),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_3982),
.B(n_163),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_3954),
.Y(n_4211)
);

BUFx2_ASAP7_75t_L g4212 ( 
.A(n_3997),
.Y(n_4212)
);

AOI22xp33_ASAP7_75t_L g4213 ( 
.A1(n_3940),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3937),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3937),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_3946),
.B(n_165),
.Y(n_4216)
);

OAI22xp33_ASAP7_75t_L g4217 ( 
.A1(n_4152),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_4217)
);

OAI221xp5_ASAP7_75t_L g4218 ( 
.A1(n_4188),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_4218)
);

BUFx2_ASAP7_75t_L g4219 ( 
.A(n_4189),
.Y(n_4219)
);

OAI22xp5_ASAP7_75t_SL g4220 ( 
.A1(n_4141),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.Y(n_4220)
);

OAI211xp5_ASAP7_75t_L g4221 ( 
.A1(n_4131),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_4221)
);

AOI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4154),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_4222)
);

NAND4xp25_ASAP7_75t_L g4223 ( 
.A(n_4092),
.B(n_180),
.C(n_181),
.D(n_179),
.Y(n_4223)
);

AOI22xp33_ASAP7_75t_L g4224 ( 
.A1(n_4137),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_4224)
);

AOI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_4140),
.A2(n_182),
.B1(n_178),
.B2(n_181),
.Y(n_4225)
);

AOI211xp5_ASAP7_75t_SL g4226 ( 
.A1(n_4208),
.A2(n_186),
.B(n_182),
.C(n_185),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_4175),
.Y(n_4227)
);

OAI211xp5_ASAP7_75t_L g4228 ( 
.A1(n_4213),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4193),
.B(n_187),
.Y(n_4229)
);

OAI31xp33_ASAP7_75t_SL g4230 ( 
.A1(n_4203),
.A2(n_191),
.A3(n_192),
.B(n_190),
.Y(n_4230)
);

OAI33xp33_ASAP7_75t_L g4231 ( 
.A1(n_4109),
.A2(n_4112),
.A3(n_4100),
.B1(n_4114),
.B2(n_4163),
.B3(n_4119),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4082),
.Y(n_4232)
);

INVxp67_ASAP7_75t_SL g4233 ( 
.A(n_4088),
.Y(n_4233)
);

BUFx3_ASAP7_75t_L g4234 ( 
.A(n_4202),
.Y(n_4234)
);

NOR2xp33_ASAP7_75t_R g4235 ( 
.A(n_4202),
.B(n_189),
.Y(n_4235)
);

AOI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_4168),
.A2(n_192),
.B1(n_189),
.B2(n_190),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_4120),
.B(n_193),
.Y(n_4237)
);

OAI22xp5_ASAP7_75t_SL g4238 ( 
.A1(n_4093),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_4238)
);

OAI211xp5_ASAP7_75t_L g4239 ( 
.A1(n_4159),
.A2(n_197),
.B(n_194),
.C(n_196),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4202),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4084),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4156),
.A2(n_201),
.B1(n_198),
.B2(n_200),
.Y(n_4242)
);

NAND4xp25_ASAP7_75t_L g4243 ( 
.A(n_4161),
.B(n_4136),
.C(n_4125),
.D(n_4128),
.Y(n_4243)
);

AND2x2_ASAP7_75t_SL g4244 ( 
.A(n_4145),
.B(n_200),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4101),
.Y(n_4245)
);

OAI332xp33_ASAP7_75t_L g4246 ( 
.A1(n_4165),
.A2(n_206),
.A3(n_205),
.B1(n_203),
.B2(n_207),
.B3(n_201),
.C1(n_202),
.C2(n_204),
.Y(n_4246)
);

NOR2xp33_ASAP7_75t_L g4247 ( 
.A(n_4094),
.B(n_203),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_4129),
.A2(n_204),
.B(n_205),
.Y(n_4248)
);

OAI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_4126),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_4249)
);

BUFx2_ASAP7_75t_L g4250 ( 
.A(n_4204),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4080),
.B(n_209),
.Y(n_4251)
);

OAI322xp33_ASAP7_75t_L g4252 ( 
.A1(n_4110),
.A2(n_4106),
.A3(n_4143),
.B1(n_4146),
.B2(n_4139),
.C1(n_4123),
.C2(n_4155),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4065),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_4212),
.B(n_210),
.Y(n_4254)
);

NAND3xp33_ASAP7_75t_L g4255 ( 
.A(n_4081),
.B(n_211),
.C(n_213),
.Y(n_4255)
);

NOR2xp33_ASAP7_75t_R g4256 ( 
.A(n_4172),
.B(n_211),
.Y(n_4256)
);

OAI211xp5_ASAP7_75t_L g4257 ( 
.A1(n_4102),
.A2(n_216),
.B(n_213),
.C(n_215),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4074),
.Y(n_4258)
);

AO21x2_ASAP7_75t_L g4259 ( 
.A1(n_4170),
.A2(n_215),
.B(n_217),
.Y(n_4259)
);

OAI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4121),
.A2(n_217),
.B(n_218),
.Y(n_4260)
);

AOI33xp33_ASAP7_75t_L g4261 ( 
.A1(n_4138),
.A2(n_220),
.A3(n_222),
.B1(n_218),
.B2(n_219),
.B3(n_221),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4075),
.Y(n_4262)
);

AOI31xp33_ASAP7_75t_L g4263 ( 
.A1(n_4098),
.A2(n_223),
.A3(n_220),
.B(n_222),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4077),
.Y(n_4264)
);

AOI22xp33_ASAP7_75t_L g4265 ( 
.A1(n_4158),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4078),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4057),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4085),
.Y(n_4268)
);

OR2x6_ASAP7_75t_L g4269 ( 
.A(n_4067),
.B(n_224),
.Y(n_4269)
);

OAI31xp33_ASAP7_75t_L g4270 ( 
.A1(n_4197),
.A2(n_228),
.A3(n_225),
.B(n_226),
.Y(n_4270)
);

AOI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4162),
.A2(n_230),
.B1(n_226),
.B2(n_228),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_4124),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_4272)
);

AOI211x1_ASAP7_75t_L g4273 ( 
.A1(n_4118),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4058),
.Y(n_4274)
);

NOR2x1_ASAP7_75t_SL g4275 ( 
.A(n_4073),
.B(n_235),
.Y(n_4275)
);

OAI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4127),
.A2(n_239),
.B1(n_235),
.B2(n_237),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4172),
.Y(n_4277)
);

NAND3xp33_ASAP7_75t_L g4278 ( 
.A(n_4105),
.B(n_239),
.C(n_240),
.Y(n_4278)
);

OR2x2_ASAP7_75t_L g4279 ( 
.A(n_4103),
.B(n_241),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4061),
.B(n_242),
.Y(n_4280)
);

AOI22xp33_ASAP7_75t_SL g4281 ( 
.A1(n_4068),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_4281)
);

AO21x1_ASAP7_75t_L g4282 ( 
.A1(n_4108),
.A2(n_243),
.B(n_244),
.Y(n_4282)
);

BUFx3_ASAP7_75t_L g4283 ( 
.A(n_4111),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4086),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4063),
.Y(n_4285)
);

OAI211xp5_ASAP7_75t_L g4286 ( 
.A1(n_4149),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_4286)
);

OAI22xp33_ASAP7_75t_L g4287 ( 
.A1(n_4115),
.A2(n_4113),
.B1(n_4195),
.B2(n_4079),
.Y(n_4287)
);

AOI22xp33_ASAP7_75t_SL g4288 ( 
.A1(n_4060),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_4288)
);

NAND4xp25_ASAP7_75t_L g4289 ( 
.A(n_4116),
.B(n_250),
.C(n_251),
.D(n_249),
.Y(n_4289)
);

AOI22xp33_ASAP7_75t_L g4290 ( 
.A1(n_4142),
.A2(n_252),
.B1(n_248),
.B2(n_251),
.Y(n_4290)
);

BUFx2_ASAP7_75t_L g4291 ( 
.A(n_4097),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4089),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4099),
.Y(n_4293)
);

AND2x4_ASAP7_75t_L g4294 ( 
.A(n_4062),
.B(n_252),
.Y(n_4294)
);

INVxp67_ASAP7_75t_SL g4295 ( 
.A(n_4091),
.Y(n_4295)
);

OAI22xp5_ASAP7_75t_SL g4296 ( 
.A1(n_4132),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_4296)
);

INVxp67_ASAP7_75t_L g4297 ( 
.A(n_4072),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4171),
.Y(n_4298)
);

HB1xp67_ASAP7_75t_L g4299 ( 
.A(n_4090),
.Y(n_4299)
);

NOR2x1_ASAP7_75t_L g4300 ( 
.A(n_4056),
.B(n_253),
.Y(n_4300)
);

AOI22xp33_ASAP7_75t_SL g4301 ( 
.A1(n_4150),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_4301)
);

AOI22xp33_ASAP7_75t_L g4302 ( 
.A1(n_4135),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4182),
.Y(n_4303)
);

NAND3xp33_ASAP7_75t_L g4304 ( 
.A(n_4122),
.B(n_258),
.C(n_259),
.Y(n_4304)
);

AOI22xp33_ASAP7_75t_L g4305 ( 
.A1(n_4133),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4184),
.Y(n_4306)
);

INVx4_ASAP7_75t_SL g4307 ( 
.A(n_4070),
.Y(n_4307)
);

AOI22xp33_ASAP7_75t_L g4308 ( 
.A1(n_4153),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4308)
);

OR2x2_ASAP7_75t_L g4309 ( 
.A(n_4064),
.B(n_264),
.Y(n_4309)
);

NOR2xp67_ASAP7_75t_L g4310 ( 
.A(n_4185),
.B(n_265),
.Y(n_4310)
);

OAI22xp5_ASAP7_75t_L g4311 ( 
.A1(n_4173),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_4311)
);

INVxp67_ASAP7_75t_SL g4312 ( 
.A(n_4083),
.Y(n_4312)
);

AOI22xp33_ASAP7_75t_L g4313 ( 
.A1(n_4157),
.A2(n_4167),
.B1(n_4151),
.B2(n_4130),
.Y(n_4313)
);

OR2x6_ASAP7_75t_L g4314 ( 
.A(n_4055),
.B(n_266),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4087),
.Y(n_4315)
);

NOR2xp33_ASAP7_75t_L g4316 ( 
.A(n_4104),
.B(n_267),
.Y(n_4316)
);

INVx1_ASAP7_75t_SL g4317 ( 
.A(n_4176),
.Y(n_4317)
);

OR2x2_ASAP7_75t_L g4318 ( 
.A(n_4169),
.B(n_268),
.Y(n_4318)
);

AOI221xp5_ASAP7_75t_L g4319 ( 
.A1(n_4148),
.A2(n_272),
.B1(n_269),
.B2(n_271),
.C(n_273),
.Y(n_4319)
);

AO21x2_ASAP7_75t_L g4320 ( 
.A1(n_4174),
.A2(n_269),
.B(n_271),
.Y(n_4320)
);

NOR2x1_ASAP7_75t_L g4321 ( 
.A(n_4196),
.B(n_273),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4187),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4190),
.Y(n_4323)
);

INVx1_ASAP7_75t_SL g4324 ( 
.A(n_4179),
.Y(n_4324)
);

OA21x2_ASAP7_75t_L g4325 ( 
.A1(n_4191),
.A2(n_274),
.B(n_275),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_4160),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4211),
.Y(n_4327)
);

AOI22xp33_ASAP7_75t_L g4328 ( 
.A1(n_4147),
.A2(n_4134),
.B1(n_4144),
.B2(n_4164),
.Y(n_4328)
);

NAND3xp33_ASAP7_75t_SL g4329 ( 
.A(n_4069),
.B(n_276),
.C(n_277),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4194),
.Y(n_4330)
);

OAI211xp5_ASAP7_75t_L g4331 ( 
.A1(n_4177),
.A2(n_280),
.B(n_277),
.C(n_278),
.Y(n_4331)
);

AOI22xp33_ASAP7_75t_L g4332 ( 
.A1(n_4166),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4332)
);

OAI22xp5_ASAP7_75t_L g4333 ( 
.A1(n_4178),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_4333)
);

NAND3xp33_ASAP7_75t_L g4334 ( 
.A(n_4216),
.B(n_4183),
.C(n_4180),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4096),
.B(n_283),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4199),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4181),
.B(n_284),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_4059),
.B(n_285),
.Y(n_4338)
);

AND2x4_ASAP7_75t_L g4339 ( 
.A(n_4192),
.B(n_285),
.Y(n_4339)
);

AND2x2_ASAP7_75t_L g4340 ( 
.A(n_4210),
.B(n_286),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4071),
.B(n_286),
.Y(n_4341)
);

AOI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4200),
.A2(n_290),
.B1(n_287),
.B2(n_289),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4076),
.B(n_289),
.Y(n_4343)
);

OAI221xp5_ASAP7_75t_L g4344 ( 
.A1(n_4107),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.C(n_294),
.Y(n_4344)
);

BUFx6f_ASAP7_75t_L g4345 ( 
.A(n_4186),
.Y(n_4345)
);

OAI22xp33_ASAP7_75t_L g4346 ( 
.A1(n_4198),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_R g4347 ( 
.A(n_4095),
.B(n_296),
.Y(n_4347)
);

INVxp67_ASAP7_75t_SL g4348 ( 
.A(n_4205),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4206),
.A2(n_297),
.B(n_298),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_4209),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4214),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4215),
.B(n_297),
.Y(n_4352)
);

INVx2_ASAP7_75t_SL g4353 ( 
.A(n_4117),
.Y(n_4353)
);

AOI21x1_ASAP7_75t_L g4354 ( 
.A1(n_4201),
.A2(n_298),
.B(n_300),
.Y(n_4354)
);

INVx2_ASAP7_75t_SL g4355 ( 
.A(n_4066),
.Y(n_4355)
);

AOI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4207),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_4356)
);

NAND3xp33_ASAP7_75t_L g4357 ( 
.A(n_4188),
.B(n_301),
.C(n_304),
.Y(n_4357)
);

OAI211xp5_ASAP7_75t_L g4358 ( 
.A1(n_4188),
.A2(n_306),
.B(n_304),
.C(n_305),
.Y(n_4358)
);

OAI332xp33_ASAP7_75t_L g4359 ( 
.A1(n_4152),
.A2(n_311),
.A3(n_310),
.B1(n_308),
.B2(n_312),
.B3(n_305),
.C1(n_307),
.C2(n_309),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4082),
.Y(n_4360)
);

AND2x4_ASAP7_75t_L g4361 ( 
.A(n_4120),
.B(n_307),
.Y(n_4361)
);

NOR2x1_ASAP7_75t_R g4362 ( 
.A(n_4202),
.B(n_308),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4140),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4189),
.B(n_309),
.Y(n_4364)
);

BUFx3_ASAP7_75t_L g4365 ( 
.A(n_4202),
.Y(n_4365)
);

AND2x2_ASAP7_75t_SL g4366 ( 
.A(n_4131),
.B(n_310),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_4175),
.Y(n_4367)
);

INVxp67_ASAP7_75t_L g4368 ( 
.A(n_4140),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4082),
.Y(n_4369)
);

OAI221xp5_ASAP7_75t_L g4370 ( 
.A1(n_4188),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.C(n_314),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4082),
.Y(n_4371)
);

BUFx2_ASAP7_75t_L g4372 ( 
.A(n_4189),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4202),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4131),
.B(n_314),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4082),
.Y(n_4375)
);

INVx2_ASAP7_75t_SL g4376 ( 
.A(n_4202),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4202),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4202),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4082),
.Y(n_4379)
);

BUFx2_ASAP7_75t_L g4380 ( 
.A(n_4189),
.Y(n_4380)
);

HB1xp67_ASAP7_75t_L g4381 ( 
.A(n_4175),
.Y(n_4381)
);

NAND2x1_ASAP7_75t_L g4382 ( 
.A(n_4189),
.B(n_315),
.Y(n_4382)
);

OAI332xp33_ASAP7_75t_L g4383 ( 
.A1(n_4152),
.A2(n_323),
.A3(n_322),
.B1(n_319),
.B2(n_324),
.B3(n_316),
.C1(n_317),
.C2(n_320),
.Y(n_4383)
);

INVxp67_ASAP7_75t_L g4384 ( 
.A(n_4140),
.Y(n_4384)
);

OAI31xp33_ASAP7_75t_L g4385 ( 
.A1(n_4188),
.A2(n_320),
.A3(n_316),
.B(n_319),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4082),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4152),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4131),
.B(n_325),
.Y(n_4388)
);

OAI211xp5_ASAP7_75t_L g4389 ( 
.A1(n_4188),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_4389)
);

OR2x6_ASAP7_75t_L g4390 ( 
.A(n_4140),
.B(n_327),
.Y(n_4390)
);

AOI322xp5_ASAP7_75t_L g4391 ( 
.A1(n_4152),
.A2(n_333),
.A3(n_332),
.B1(n_330),
.B2(n_328),
.C1(n_329),
.C2(n_331),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4131),
.B(n_328),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4202),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4131),
.B(n_330),
.Y(n_4394)
);

BUFx8_ASAP7_75t_L g4395 ( 
.A(n_4116),
.Y(n_4395)
);

INVx2_ASAP7_75t_SL g4396 ( 
.A(n_4202),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_4152),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4131),
.B(n_335),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4189),
.B(n_335),
.Y(n_4399)
);

OR2x2_ASAP7_75t_L g4400 ( 
.A(n_4080),
.B(n_336),
.Y(n_4400)
);

NAND4xp25_ASAP7_75t_SL g4401 ( 
.A(n_4092),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_R g4402 ( 
.A(n_4202),
.B(n_337),
.Y(n_4402)
);

OAI22xp5_ASAP7_75t_L g4403 ( 
.A1(n_4152),
.A2(n_341),
.B1(n_338),
.B2(n_340),
.Y(n_4403)
);

BUFx3_ASAP7_75t_L g4404 ( 
.A(n_4202),
.Y(n_4404)
);

OAI33xp33_ASAP7_75t_L g4405 ( 
.A1(n_4208),
.A2(n_345),
.A3(n_347),
.B1(n_342),
.B2(n_344),
.B3(n_346),
.Y(n_4405)
);

BUFx3_ASAP7_75t_L g4406 ( 
.A(n_4202),
.Y(n_4406)
);

HB1xp67_ASAP7_75t_L g4407 ( 
.A(n_4175),
.Y(n_4407)
);

NOR2xp67_ASAP7_75t_L g4408 ( 
.A(n_4202),
.B(n_342),
.Y(n_4408)
);

OAI221xp5_ASAP7_75t_L g4409 ( 
.A1(n_4188),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.C(n_347),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4131),
.B(n_348),
.Y(n_4410)
);

INVx3_ASAP7_75t_SL g4411 ( 
.A(n_4202),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_4283),
.B(n_348),
.Y(n_4412)
);

AOI21x1_ASAP7_75t_L g4413 ( 
.A1(n_4390),
.A2(n_357),
.B(n_349),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4307),
.B(n_349),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4231),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_4415)
);

HB1xp67_ASAP7_75t_L g4416 ( 
.A(n_4219),
.Y(n_4416)
);

NOR3xp33_ASAP7_75t_L g4417 ( 
.A(n_4246),
.B(n_350),
.C(n_353),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4234),
.Y(n_4418)
);

OAI211xp5_ASAP7_75t_SL g4419 ( 
.A1(n_4230),
.A2(n_355),
.B(n_353),
.C(n_354),
.Y(n_4419)
);

NAND3xp33_ASAP7_75t_L g4420 ( 
.A(n_4226),
.B(n_4385),
.C(n_4391),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4250),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4243),
.A2(n_358),
.B1(n_354),
.B2(n_356),
.Y(n_4422)
);

NAND3xp33_ASAP7_75t_L g4423 ( 
.A(n_4255),
.B(n_356),
.C(n_358),
.Y(n_4423)
);

AND2x4_ASAP7_75t_L g4424 ( 
.A(n_4365),
.B(n_359),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4307),
.B(n_359),
.Y(n_4425)
);

NOR3xp33_ASAP7_75t_L g4426 ( 
.A(n_4252),
.B(n_360),
.C(n_361),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_L g4427 ( 
.A(n_4411),
.B(n_361),
.Y(n_4427)
);

AOI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_4363),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_4428)
);

NAND4xp75_ASAP7_75t_L g4429 ( 
.A(n_4282),
.B(n_368),
.C(n_365),
.D(n_366),
.Y(n_4429)
);

NAND4xp75_ASAP7_75t_L g4430 ( 
.A(n_4366),
.B(n_369),
.C(n_366),
.D(n_368),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4368),
.B(n_369),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4233),
.B(n_370),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4404),
.Y(n_4433)
);

OR2x2_ASAP7_75t_L g4434 ( 
.A(n_4295),
.B(n_4291),
.Y(n_4434)
);

NOR3xp33_ASAP7_75t_SL g4435 ( 
.A(n_4287),
.B(n_370),
.C(n_372),
.Y(n_4435)
);

NOR2x1_ASAP7_75t_L g4436 ( 
.A(n_4390),
.B(n_373),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4227),
.Y(n_4437)
);

NOR3xp33_ASAP7_75t_L g4438 ( 
.A(n_4359),
.B(n_373),
.C(n_374),
.Y(n_4438)
);

AND2x4_ASAP7_75t_L g4439 ( 
.A(n_4406),
.B(n_374),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4367),
.Y(n_4440)
);

AOI22xp33_ASAP7_75t_SL g4441 ( 
.A1(n_4244),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4441)
);

OR2x2_ASAP7_75t_SL g4442 ( 
.A(n_4357),
.B(n_376),
.Y(n_4442)
);

NOR2xp33_ASAP7_75t_L g4443 ( 
.A(n_4345),
.B(n_377),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4372),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4381),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4384),
.B(n_379),
.Y(n_4446)
);

NAND4xp25_ASAP7_75t_L g4447 ( 
.A(n_4387),
.B(n_381),
.C(n_379),
.D(n_380),
.Y(n_4447)
);

AOI221xp5_ASAP7_75t_L g4448 ( 
.A1(n_4220),
.A2(n_383),
.B1(n_380),
.B2(n_382),
.C(n_384),
.Y(n_4448)
);

OAI211xp5_ASAP7_75t_SL g4449 ( 
.A1(n_4328),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_4449)
);

INVx5_ASAP7_75t_L g4450 ( 
.A(n_4376),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4407),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_L g4452 ( 
.A1(n_4267),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4452)
);

AO21x2_ASAP7_75t_L g4453 ( 
.A1(n_4374),
.A2(n_386),
.B(n_388),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4324),
.B(n_388),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4380),
.B(n_389),
.Y(n_4455)
);

AOI22xp5_ASAP7_75t_L g4456 ( 
.A1(n_4238),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4240),
.B(n_392),
.Y(n_4457)
);

INVx3_ASAP7_75t_L g4458 ( 
.A(n_4345),
.Y(n_4458)
);

NAND4xp75_ASAP7_75t_L g4459 ( 
.A(n_4273),
.B(n_395),
.C(n_393),
.D(n_394),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4373),
.B(n_393),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4377),
.B(n_394),
.Y(n_4461)
);

NAND4xp75_ASAP7_75t_L g4462 ( 
.A(n_4225),
.B(n_401),
.C(n_396),
.D(n_398),
.Y(n_4462)
);

OAI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_4218),
.A2(n_403),
.B1(n_398),
.B2(n_402),
.Y(n_4463)
);

OAI211xp5_ASAP7_75t_SL g4464 ( 
.A1(n_4260),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4378),
.B(n_405),
.Y(n_4465)
);

AOI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_4396),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4466)
);

AOI22xp33_ASAP7_75t_L g4467 ( 
.A1(n_4274),
.A2(n_411),
.B1(n_408),
.B2(n_410),
.Y(n_4467)
);

NAND3xp33_ASAP7_75t_L g4468 ( 
.A(n_4319),
.B(n_410),
.C(n_411),
.Y(n_4468)
);

AOI22xp33_ASAP7_75t_L g4469 ( 
.A1(n_4278),
.A2(n_4405),
.B1(n_4223),
.B2(n_4401),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4355),
.B(n_412),
.Y(n_4470)
);

NAND3xp33_ASAP7_75t_L g4471 ( 
.A(n_4239),
.B(n_4221),
.C(n_4358),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4312),
.B(n_412),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4259),
.B(n_413),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4393),
.Y(n_4474)
);

AOI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_4296),
.A2(n_4389),
.B1(n_4257),
.B2(n_4370),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4277),
.B(n_4348),
.Y(n_4476)
);

OR2x2_ASAP7_75t_L g4477 ( 
.A(n_4297),
.B(n_413),
.Y(n_4477)
);

OR2x2_ASAP7_75t_L g4478 ( 
.A(n_4251),
.B(n_414),
.Y(n_4478)
);

OAI211xp5_ASAP7_75t_L g4479 ( 
.A1(n_4270),
.A2(n_4402),
.B(n_4235),
.C(n_4222),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4353),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4229),
.B(n_415),
.Y(n_4481)
);

NAND2xp33_ASAP7_75t_SL g4482 ( 
.A(n_4382),
.B(n_415),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4254),
.B(n_417),
.Y(n_4483)
);

BUFx3_ASAP7_75t_L g4484 ( 
.A(n_4395),
.Y(n_4484)
);

NAND3xp33_ASAP7_75t_L g4485 ( 
.A(n_4261),
.B(n_418),
.C(n_419),
.Y(n_4485)
);

AOI22x1_ASAP7_75t_L g4486 ( 
.A1(n_4248),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_4486)
);

AOI22xp33_ASAP7_75t_SL g4487 ( 
.A1(n_4409),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4320),
.B(n_421),
.Y(n_4488)
);

AO21x2_ASAP7_75t_L g4489 ( 
.A1(n_4388),
.A2(n_423),
.B(n_424),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4280),
.Y(n_4490)
);

NAND3xp33_ASAP7_75t_SL g4491 ( 
.A(n_4349),
.B(n_424),
.C(n_425),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4364),
.B(n_425),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4350),
.Y(n_4493)
);

AOI211xp5_ASAP7_75t_L g4494 ( 
.A1(n_4383),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4310),
.B(n_426),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4253),
.Y(n_4496)
);

OAI221xp5_ASAP7_75t_L g4497 ( 
.A1(n_4344),
.A2(n_433),
.B1(n_430),
.B2(n_431),
.C(n_434),
.Y(n_4497)
);

NAND3xp33_ASAP7_75t_SL g4498 ( 
.A(n_4286),
.B(n_431),
.C(n_433),
.Y(n_4498)
);

AOI22xp33_ASAP7_75t_L g4499 ( 
.A1(n_4304),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_4275),
.B(n_435),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4258),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4392),
.B(n_436),
.Y(n_4502)
);

NAND4xp75_ASAP7_75t_L g4503 ( 
.A(n_4408),
.B(n_439),
.C(n_437),
.D(n_438),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4262),
.Y(n_4504)
);

OAI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_4241),
.A2(n_438),
.B(n_439),
.Y(n_4505)
);

INVxp67_ASAP7_75t_L g4506 ( 
.A(n_4362),
.Y(n_4506)
);

NAND4xp75_ASAP7_75t_L g4507 ( 
.A(n_4300),
.B(n_444),
.C(n_440),
.D(n_442),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4399),
.B(n_440),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4317),
.B(n_442),
.Y(n_4509)
);

OAI21xp5_ASAP7_75t_L g4510 ( 
.A1(n_4263),
.A2(n_4321),
.B(n_4394),
.Y(n_4510)
);

NAND3xp33_ASAP7_75t_L g4511 ( 
.A(n_4281),
.B(n_444),
.C(n_445),
.Y(n_4511)
);

AOI22xp33_ASAP7_75t_L g4512 ( 
.A1(n_4334),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_4512)
);

NAND3xp33_ASAP7_75t_L g4513 ( 
.A(n_4228),
.B(n_446),
.C(n_447),
.Y(n_4513)
);

AND2x4_ASAP7_75t_L g4514 ( 
.A(n_4232),
.B(n_448),
.Y(n_4514)
);

OR2x2_ASAP7_75t_L g4515 ( 
.A(n_4400),
.B(n_448),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4299),
.B(n_4285),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_4237),
.Y(n_4517)
);

NAND4xp25_ASAP7_75t_SL g4518 ( 
.A(n_4397),
.B(n_451),
.C(n_449),
.D(n_450),
.Y(n_4518)
);

OAI211xp5_ASAP7_75t_SL g4519 ( 
.A1(n_4313),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4315),
.B(n_452),
.Y(n_4520)
);

NOR3xp33_ASAP7_75t_L g4521 ( 
.A(n_4331),
.B(n_4329),
.C(n_4289),
.Y(n_4521)
);

OA211x2_ASAP7_75t_L g4522 ( 
.A1(n_4398),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_4522)
);

NAND3xp33_ASAP7_75t_L g4523 ( 
.A(n_4242),
.B(n_453),
.C(n_454),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4327),
.B(n_455),
.Y(n_4524)
);

NAND3xp33_ASAP7_75t_L g4525 ( 
.A(n_4224),
.B(n_456),
.C(n_457),
.Y(n_4525)
);

OR2x2_ASAP7_75t_L g4526 ( 
.A(n_4245),
.B(n_456),
.Y(n_4526)
);

OAI211xp5_ASAP7_75t_SL g4527 ( 
.A1(n_4410),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_4527)
);

AOI22xp33_ASAP7_75t_L g4528 ( 
.A1(n_4301),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_4528)
);

OAI211xp5_ASAP7_75t_L g4529 ( 
.A1(n_4288),
.A2(n_4302),
.B(n_4342),
.C(n_4308),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4341),
.B(n_464),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4352),
.B(n_464),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4337),
.B(n_4340),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4339),
.B(n_465),
.Y(n_4533)
);

AOI22xp5_ASAP7_75t_L g4534 ( 
.A1(n_4217),
.A2(n_469),
.B1(n_466),
.B2(n_467),
.Y(n_4534)
);

NAND3xp33_ASAP7_75t_SL g4535 ( 
.A(n_4347),
.B(n_467),
.C(n_469),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_4360),
.B(n_470),
.Y(n_4536)
);

AOI22xp33_ASAP7_75t_L g4537 ( 
.A1(n_4311),
.A2(n_473),
.B1(n_470),
.B2(n_472),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4369),
.B(n_472),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4371),
.B(n_474),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_SL g4540 ( 
.A(n_4346),
.B(n_475),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4375),
.B(n_475),
.Y(n_4541)
);

OAI211xp5_ASAP7_75t_SL g4542 ( 
.A1(n_4326),
.A2(n_478),
.B(n_476),
.C(n_477),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4333),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_4543)
);

OR2x2_ASAP7_75t_L g4544 ( 
.A(n_4379),
.B(n_480),
.Y(n_4544)
);

AOI22xp33_ASAP7_75t_SL g4545 ( 
.A1(n_4325),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_4545)
);

OR2x2_ASAP7_75t_L g4546 ( 
.A(n_4386),
.B(n_4279),
.Y(n_4546)
);

OAI211xp5_ASAP7_75t_SL g4547 ( 
.A1(n_4356),
.A2(n_485),
.B(n_482),
.C(n_484),
.Y(n_4547)
);

OR2x2_ASAP7_75t_L g4548 ( 
.A(n_4309),
.B(n_486),
.Y(n_4548)
);

OR2x2_ASAP7_75t_L g4549 ( 
.A(n_4434),
.B(n_4318),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4484),
.B(n_4269),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4458),
.B(n_4269),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4416),
.B(n_4421),
.Y(n_4552)
);

OR2x2_ASAP7_75t_L g4553 ( 
.A(n_4444),
.B(n_4264),
.Y(n_4553)
);

INVx8_ASAP7_75t_L g4554 ( 
.A(n_4424),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4517),
.B(n_4314),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4437),
.B(n_4266),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_4450),
.Y(n_4557)
);

INVx1_ASAP7_75t_SL g4558 ( 
.A(n_4482),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4440),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4415),
.B(n_4316),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4532),
.B(n_4314),
.Y(n_4561)
);

OAI211xp5_ASAP7_75t_SL g4562 ( 
.A1(n_4494),
.A2(n_4290),
.B(n_4265),
.C(n_4343),
.Y(n_4562)
);

NAND3xp33_ASAP7_75t_L g4563 ( 
.A(n_4426),
.B(n_4271),
.C(n_4236),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4445),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4451),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4536),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4418),
.B(n_4247),
.Y(n_4567)
);

NOR3xp33_ASAP7_75t_L g4568 ( 
.A(n_4417),
.B(n_4249),
.C(n_4272),
.Y(n_4568)
);

HB1xp67_ASAP7_75t_L g4569 ( 
.A(n_4450),
.Y(n_4569)
);

BUFx3_ASAP7_75t_L g4570 ( 
.A(n_4450),
.Y(n_4570)
);

INVx3_ASAP7_75t_L g4571 ( 
.A(n_4433),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4480),
.Y(n_4572)
);

AND2x4_ASAP7_75t_L g4573 ( 
.A(n_4506),
.B(n_4361),
.Y(n_4573)
);

BUFx2_ASAP7_75t_L g4574 ( 
.A(n_4436),
.Y(n_4574)
);

AOI222xp33_ASAP7_75t_L g4575 ( 
.A1(n_4420),
.A2(n_4403),
.B1(n_4276),
.B2(n_4305),
.C1(n_4332),
.C2(n_4335),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4539),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4541),
.Y(n_4577)
);

OAI211xp5_ASAP7_75t_L g4578 ( 
.A1(n_4438),
.A2(n_4256),
.B(n_4325),
.C(n_4354),
.Y(n_4578)
);

HB1xp67_ASAP7_75t_L g4579 ( 
.A(n_4414),
.Y(n_4579)
);

BUFx2_ASAP7_75t_L g4580 ( 
.A(n_4425),
.Y(n_4580)
);

INVx4_ASAP7_75t_L g4581 ( 
.A(n_4424),
.Y(n_4581)
);

OAI221xp5_ASAP7_75t_L g4582 ( 
.A1(n_4435),
.A2(n_4292),
.B1(n_4293),
.B2(n_4284),
.C(n_4268),
.Y(n_4582)
);

OR2x2_ASAP7_75t_L g4583 ( 
.A(n_4546),
.B(n_4298),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4476),
.B(n_4490),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4470),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4526),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4544),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4521),
.B(n_4303),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4474),
.B(n_4306),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4457),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4493),
.Y(n_4591)
);

INVx1_ASAP7_75t_SL g4592 ( 
.A(n_4455),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4510),
.B(n_4294),
.Y(n_4593)
);

OR2x2_ASAP7_75t_L g4594 ( 
.A(n_4432),
.B(n_4322),
.Y(n_4594)
);

OAI211xp5_ASAP7_75t_L g4595 ( 
.A1(n_4479),
.A2(n_4330),
.B(n_4336),
.C(n_4323),
.Y(n_4595)
);

AND2x4_ASAP7_75t_L g4596 ( 
.A(n_4460),
.B(n_4461),
.Y(n_4596)
);

OR2x2_ASAP7_75t_L g4597 ( 
.A(n_4453),
.B(n_4351),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4489),
.B(n_4338),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4477),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4520),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4431),
.B(n_486),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4524),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4446),
.B(n_4427),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4465),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4509),
.B(n_487),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4496),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4516),
.B(n_487),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4530),
.B(n_488),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4501),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4504),
.Y(n_4610)
);

HB1xp67_ASAP7_75t_L g4611 ( 
.A(n_4413),
.Y(n_4611)
);

OAI21xp5_ASAP7_75t_L g4612 ( 
.A1(n_4468),
.A2(n_488),
.B(n_489),
.Y(n_4612)
);

INVx4_ASAP7_75t_L g4613 ( 
.A(n_4439),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_SL g4614 ( 
.A(n_4430),
.B(n_490),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4514),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4548),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4481),
.B(n_490),
.Y(n_4617)
);

AND2x4_ASAP7_75t_SL g4618 ( 
.A(n_4439),
.B(n_491),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_4472),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4514),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4478),
.Y(n_4621)
);

HB1xp67_ASAP7_75t_L g4622 ( 
.A(n_4454),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4515),
.Y(n_4623)
);

AND2x4_ASAP7_75t_L g4624 ( 
.A(n_4533),
.B(n_491),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4483),
.B(n_492),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4492),
.B(n_493),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4538),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_L g4628 ( 
.A(n_4469),
.B(n_494),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4531),
.Y(n_4629)
);

INVx3_ASAP7_75t_L g4630 ( 
.A(n_4508),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4473),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4412),
.B(n_495),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4488),
.Y(n_4633)
);

OAI21xp33_ASAP7_75t_L g4634 ( 
.A1(n_4475),
.A2(n_495),
.B(n_496),
.Y(n_4634)
);

NOR3xp33_ASAP7_75t_L g4635 ( 
.A(n_4498),
.B(n_496),
.C(n_497),
.Y(n_4635)
);

INVx2_ASAP7_75t_SL g4636 ( 
.A(n_4500),
.Y(n_4636)
);

HB1xp67_ASAP7_75t_L g4637 ( 
.A(n_4429),
.Y(n_4637)
);

AOI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4419),
.A2(n_500),
.B1(n_497),
.B2(n_499),
.Y(n_4638)
);

OAI221xp5_ASAP7_75t_L g4639 ( 
.A1(n_4529),
.A2(n_502),
.B1(n_499),
.B2(n_500),
.C(n_503),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4502),
.Y(n_4640)
);

AND2x4_ASAP7_75t_L g4641 ( 
.A(n_4443),
.B(n_502),
.Y(n_4641)
);

OAI21xp33_ASAP7_75t_SL g4642 ( 
.A1(n_4611),
.A2(n_4597),
.B(n_4558),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4620),
.Y(n_4643)
);

BUFx3_ASAP7_75t_L g4644 ( 
.A(n_4554),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4580),
.B(n_4422),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4550),
.B(n_4540),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4574),
.B(n_4471),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4573),
.B(n_4495),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4570),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4569),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4579),
.B(n_4592),
.Y(n_4651)
);

NAND5xp2_ASAP7_75t_L g4652 ( 
.A(n_4584),
.B(n_4487),
.C(n_4441),
.D(n_4448),
.E(n_4528),
.Y(n_4652)
);

XOR2x2_ASAP7_75t_L g4653 ( 
.A(n_4568),
.B(n_4485),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4637),
.B(n_4428),
.Y(n_4654)
);

INVx5_ASAP7_75t_L g4655 ( 
.A(n_4557),
.Y(n_4655)
);

OAI22xp5_ASAP7_75t_L g4656 ( 
.A1(n_4563),
.A2(n_4545),
.B1(n_4511),
.B2(n_4513),
.Y(n_4656)
);

INVx2_ASAP7_75t_SL g4657 ( 
.A(n_4554),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4581),
.B(n_4535),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4552),
.Y(n_4659)
);

INVx2_ASAP7_75t_SL g4660 ( 
.A(n_4618),
.Y(n_4660)
);

O2A1O1Ixp5_ASAP7_75t_R g4661 ( 
.A1(n_4588),
.A2(n_4442),
.B(n_4518),
.C(n_4459),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4615),
.B(n_4456),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4566),
.Y(n_4663)
);

OA222x2_ASAP7_75t_L g4664 ( 
.A1(n_4598),
.A2(n_4527),
.B1(n_4522),
.B2(n_4507),
.C1(n_4503),
.C2(n_4491),
.Y(n_4664)
);

NAND2x2_ASAP7_75t_L g4665 ( 
.A(n_4636),
.B(n_4447),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_SL g4666 ( 
.A(n_4613),
.B(n_4423),
.Y(n_4666)
);

XNOR2x1_ASAP7_75t_L g4667 ( 
.A(n_4612),
.B(n_4462),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4576),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4577),
.Y(n_4669)
);

INVxp67_ASAP7_75t_L g4670 ( 
.A(n_4614),
.Y(n_4670)
);

INVxp67_ASAP7_75t_L g4671 ( 
.A(n_4551),
.Y(n_4671)
);

AOI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4578),
.A2(n_4464),
.B1(n_4519),
.B2(n_4449),
.Y(n_4672)
);

INVxp67_ASAP7_75t_L g4673 ( 
.A(n_4561),
.Y(n_4673)
);

OAI22xp33_ASAP7_75t_L g4674 ( 
.A1(n_4638),
.A2(n_4497),
.B1(n_4534),
.B2(n_4523),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4634),
.B(n_4466),
.Y(n_4675)
);

OR2x2_ASAP7_75t_L g4676 ( 
.A(n_4549),
.B(n_4505),
.Y(n_4676)
);

INVx3_ASAP7_75t_L g4677 ( 
.A(n_4571),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4621),
.Y(n_4678)
);

OAI33xp33_ASAP7_75t_L g4679 ( 
.A1(n_4559),
.A2(n_4564),
.A3(n_4565),
.B1(n_4591),
.B2(n_4633),
.B3(n_4631),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4616),
.Y(n_4680)
);

INVx1_ASAP7_75t_SL g4681 ( 
.A(n_4555),
.Y(n_4681)
);

INVxp67_ASAP7_75t_L g4682 ( 
.A(n_4593),
.Y(n_4682)
);

AOI22xp33_ASAP7_75t_L g4683 ( 
.A1(n_4562),
.A2(n_4547),
.B1(n_4542),
.B2(n_4525),
.Y(n_4683)
);

NOR2xp33_ASAP7_75t_L g4684 ( 
.A(n_4639),
.B(n_4463),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4630),
.B(n_4512),
.Y(n_4685)
);

INVx2_ASAP7_75t_SL g4686 ( 
.A(n_4596),
.Y(n_4686)
);

OR2x6_ASAP7_75t_L g4687 ( 
.A(n_4607),
.B(n_4486),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4583),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4623),
.Y(n_4689)
);

OAI32xp33_ASAP7_75t_L g4690 ( 
.A1(n_4635),
.A2(n_4499),
.A3(n_4543),
.B1(n_4537),
.B2(n_4452),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4567),
.B(n_4467),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4586),
.Y(n_4692)
);

OAI22xp33_ASAP7_75t_L g4693 ( 
.A1(n_4560),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4590),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4604),
.B(n_505),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_R g4696 ( 
.A(n_4603),
.B(n_506),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4587),
.Y(n_4697)
);

OAI322xp33_ASAP7_75t_L g4698 ( 
.A1(n_4628),
.A2(n_512),
.A3(n_511),
.B1(n_509),
.B2(n_507),
.C1(n_508),
.C2(n_510),
.Y(n_4698)
);

OAI33xp33_ASAP7_75t_L g4699 ( 
.A1(n_4589),
.A2(n_512),
.A3(n_515),
.B1(n_509),
.B2(n_510),
.B3(n_514),
.Y(n_4699)
);

OA222x2_ASAP7_75t_L g4700 ( 
.A1(n_4556),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.C1(n_516),
.C2(n_518),
.Y(n_4700)
);

OR2x2_ASAP7_75t_L g4701 ( 
.A(n_4572),
.B(n_515),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4600),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4646),
.B(n_4622),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4660),
.B(n_4575),
.Y(n_4704)
);

INVxp67_ASAP7_75t_SL g4705 ( 
.A(n_4650),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4643),
.Y(n_4706)
);

NOR2xp67_ASAP7_75t_L g4707 ( 
.A(n_4655),
.B(n_4595),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4686),
.B(n_4602),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4681),
.B(n_4599),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4651),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4647),
.B(n_4553),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4701),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4644),
.B(n_4619),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4688),
.Y(n_4714)
);

OAI21x1_ASAP7_75t_SL g4715 ( 
.A1(n_4661),
.A2(n_4601),
.B(n_4606),
.Y(n_4715)
);

NAND2xp33_ASAP7_75t_R g4716 ( 
.A(n_4677),
.B(n_4648),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4657),
.B(n_4629),
.Y(n_4717)
);

NOR3xp33_ASAP7_75t_SL g4718 ( 
.A(n_4642),
.B(n_4627),
.C(n_4640),
.Y(n_4718)
);

NOR2xp33_ASAP7_75t_L g4719 ( 
.A(n_4670),
.B(n_4594),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4649),
.B(n_4585),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4658),
.B(n_4605),
.Y(n_4721)
);

OR2x2_ASAP7_75t_L g4722 ( 
.A(n_4654),
.B(n_4582),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4695),
.Y(n_4723)
);

AOI22xp5_ASAP7_75t_L g4724 ( 
.A1(n_4672),
.A2(n_4609),
.B1(n_4610),
.B2(n_4641),
.Y(n_4724)
);

INVx1_ASAP7_75t_SL g4725 ( 
.A(n_4655),
.Y(n_4725)
);

NOR2xp33_ASAP7_75t_L g4726 ( 
.A(n_4671),
.B(n_4617),
.Y(n_4726)
);

NOR3xp33_ASAP7_75t_L g4727 ( 
.A(n_4682),
.B(n_4632),
.C(n_4626),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4673),
.B(n_4625),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4655),
.Y(n_4729)
);

INVx1_ASAP7_75t_SL g4730 ( 
.A(n_4687),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4687),
.B(n_4608),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4689),
.Y(n_4732)
);

AOI21xp33_ASAP7_75t_SL g4733 ( 
.A1(n_4656),
.A2(n_4624),
.B(n_516),
.Y(n_4733)
);

AND2x2_ASAP7_75t_SL g4734 ( 
.A(n_4683),
.B(n_517),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4678),
.Y(n_4735)
);

NOR2xp67_ASAP7_75t_SL g4736 ( 
.A(n_4659),
.B(n_518),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4684),
.B(n_519),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4694),
.B(n_520),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4680),
.Y(n_4739)
);

AOI22xp33_ASAP7_75t_L g4740 ( 
.A1(n_4653),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4676),
.B(n_521),
.Y(n_4741)
);

AOI31xp33_ASAP7_75t_L g4742 ( 
.A1(n_4667),
.A2(n_526),
.A3(n_524),
.B(n_525),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_4652),
.B(n_524),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4692),
.Y(n_4744)
);

NOR2xp33_ASAP7_75t_L g4745 ( 
.A(n_4666),
.B(n_527),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4691),
.B(n_528),
.Y(n_4746)
);

AND2x4_ASAP7_75t_L g4747 ( 
.A(n_4697),
.B(n_529),
.Y(n_4747)
);

AOI22xp33_ASAP7_75t_L g4748 ( 
.A1(n_4665),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_4748)
);

NAND2x1p5_ASAP7_75t_L g4749 ( 
.A(n_4663),
.B(n_532),
.Y(n_4749)
);

INVx1_ASAP7_75t_SL g4750 ( 
.A(n_4725),
.Y(n_4750)
);

OR2x2_ASAP7_75t_L g4751 ( 
.A(n_4730),
.B(n_4645),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4705),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4704),
.B(n_4662),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4731),
.B(n_4675),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_SL g4755 ( 
.A(n_4707),
.B(n_4674),
.Y(n_4755)
);

AOI21xp5_ASAP7_75t_L g4756 ( 
.A1(n_4743),
.A2(n_4693),
.B(n_4690),
.Y(n_4756)
);

AOI322xp5_ASAP7_75t_L g4757 ( 
.A1(n_4718),
.A2(n_4685),
.A3(n_4702),
.B1(n_4668),
.B2(n_4669),
.C1(n_4664),
.C2(n_4700),
.Y(n_4757)
);

AOI32xp33_ASAP7_75t_L g4758 ( 
.A1(n_4748),
.A2(n_4696),
.A3(n_4679),
.B1(n_4698),
.B2(n_4699),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4728),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4729),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4703),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4709),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4708),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4713),
.B(n_532),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4734),
.B(n_533),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4726),
.B(n_4727),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4735),
.Y(n_4767)
);

HB1xp67_ASAP7_75t_L g4768 ( 
.A(n_4716),
.Y(n_4768)
);

OR2x2_ASAP7_75t_L g4769 ( 
.A(n_4722),
.B(n_4741),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_L g4770 ( 
.A(n_4733),
.B(n_533),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4711),
.B(n_534),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4717),
.B(n_534),
.Y(n_4772)
);

OR2x2_ASAP7_75t_L g4773 ( 
.A(n_4746),
.B(n_535),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4720),
.B(n_535),
.Y(n_4774)
);

OR2x2_ASAP7_75t_L g4775 ( 
.A(n_4721),
.B(n_536),
.Y(n_4775)
);

HB1xp67_ASAP7_75t_L g4776 ( 
.A(n_4749),
.Y(n_4776)
);

OR2x2_ASAP7_75t_L g4777 ( 
.A(n_4706),
.B(n_537),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4738),
.Y(n_4778)
);

OAI332xp33_ASAP7_75t_L g4779 ( 
.A1(n_4710),
.A2(n_543),
.A3(n_541),
.B1(n_539),
.B2(n_544),
.B3(n_537),
.C1(n_538),
.C2(n_540),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4719),
.B(n_538),
.Y(n_4780)
);

OR2x2_ASAP7_75t_L g4781 ( 
.A(n_4714),
.B(n_540),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4747),
.Y(n_4782)
);

NOR3xp33_ASAP7_75t_L g4783 ( 
.A(n_4712),
.B(n_543),
.C(n_544),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4742),
.B(n_545),
.Y(n_4784)
);

OR2x2_ASAP7_75t_L g4785 ( 
.A(n_4737),
.B(n_546),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4736),
.B(n_547),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4747),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4732),
.Y(n_4788)
);

AND2x2_ASAP7_75t_L g4789 ( 
.A(n_4724),
.B(n_547),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4745),
.B(n_548),
.Y(n_4790)
);

OR2x2_ASAP7_75t_L g4791 ( 
.A(n_4723),
.B(n_550),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4739),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4744),
.Y(n_4793)
);

CKINVDCx16_ASAP7_75t_R g4794 ( 
.A(n_4715),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4740),
.Y(n_4795)
);

INVx2_ASAP7_75t_SL g4796 ( 
.A(n_4729),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4705),
.B(n_550),
.Y(n_4797)
);

OAI22xp5_ASAP7_75t_L g4798 ( 
.A1(n_4794),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4755),
.A2(n_551),
.B(n_552),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4796),
.Y(n_4800)
);

AOI21xp33_ASAP7_75t_SL g4801 ( 
.A1(n_4768),
.A2(n_556),
.B(n_555),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4761),
.Y(n_4802)
);

OAI21xp33_ASAP7_75t_L g4803 ( 
.A1(n_4757),
.A2(n_554),
.B(n_557),
.Y(n_4803)
);

XNOR2x1_ASAP7_75t_L g4804 ( 
.A(n_4753),
.B(n_558),
.Y(n_4804)
);

OAI22xp5_ASAP7_75t_L g4805 ( 
.A1(n_4750),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_4805)
);

NAND3xp33_ASAP7_75t_SL g4806 ( 
.A(n_4758),
.B(n_561),
.C(n_560),
.Y(n_4806)
);

NAND2xp33_ASAP7_75t_R g4807 ( 
.A(n_4769),
.B(n_560),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4782),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4787),
.Y(n_4809)
);

AOI222xp33_ASAP7_75t_L g4810 ( 
.A1(n_4795),
.A2(n_562),
.B1(n_564),
.B2(n_559),
.C1(n_561),
.C2(n_563),
.Y(n_4810)
);

INVxp67_ASAP7_75t_L g4811 ( 
.A(n_4776),
.Y(n_4811)
);

AOI31xp33_ASAP7_75t_L g4812 ( 
.A1(n_4767),
.A2(n_565),
.A3(n_562),
.B(n_563),
.Y(n_4812)
);

OAI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_4751),
.A2(n_568),
.B1(n_565),
.B2(n_567),
.Y(n_4813)
);

NAND3xp33_ASAP7_75t_L g4814 ( 
.A(n_4756),
.B(n_4752),
.C(n_4760),
.Y(n_4814)
);

AOI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4754),
.A2(n_4766),
.B(n_4784),
.Y(n_4815)
);

AOI211xp5_ASAP7_75t_L g4816 ( 
.A1(n_4779),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4764),
.Y(n_4817)
);

OAI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4789),
.A2(n_569),
.B(n_570),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4774),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4780),
.Y(n_4820)
);

AOI211xp5_ASAP7_75t_SL g4821 ( 
.A1(n_4759),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_4821)
);

NOR2xp33_ASAP7_75t_L g4822 ( 
.A(n_4765),
.B(n_571),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4797),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4771),
.B(n_573),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4770),
.B(n_575),
.Y(n_4825)
);

AOI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4772),
.A2(n_575),
.B(n_576),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4778),
.B(n_577),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4786),
.Y(n_4828)
);

AOI31xp33_ASAP7_75t_L g4829 ( 
.A1(n_4762),
.A2(n_579),
.A3(n_577),
.B(n_578),
.Y(n_4829)
);

OAI22xp5_ASAP7_75t_L g4830 ( 
.A1(n_4763),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4781),
.Y(n_4831)
);

AOI22x1_ASAP7_75t_L g4832 ( 
.A1(n_4788),
.A2(n_4793),
.B1(n_4792),
.B2(n_4775),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4783),
.B(n_580),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4777),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4785),
.B(n_581),
.Y(n_4835)
);

AOI22xp33_ASAP7_75t_L g4836 ( 
.A1(n_4773),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4791),
.Y(n_4837)
);

NAND4xp25_ASAP7_75t_SL g4838 ( 
.A(n_4790),
.B(n_585),
.C(n_583),
.D(n_584),
.Y(n_4838)
);

NAND3xp33_ASAP7_75t_L g4839 ( 
.A(n_4757),
.B(n_584),
.C(n_585),
.Y(n_4839)
);

INVxp67_ASAP7_75t_SL g4840 ( 
.A(n_4768),
.Y(n_4840)
);

AND4x1_ASAP7_75t_L g4841 ( 
.A(n_4761),
.B(n_589),
.C(n_586),
.D(n_588),
.Y(n_4841)
);

INVxp67_ASAP7_75t_L g4842 ( 
.A(n_4768),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4750),
.B(n_586),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4761),
.Y(n_4844)
);

INVx3_ASAP7_75t_L g4845 ( 
.A(n_4782),
.Y(n_4845)
);

OAI22xp5_ASAP7_75t_L g4846 ( 
.A1(n_4794),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4761),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4761),
.Y(n_4848)
);

XNOR2x1_ASAP7_75t_L g4849 ( 
.A(n_4753),
.B(n_591),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4768),
.B(n_590),
.Y(n_4850)
);

OAI21xp33_ASAP7_75t_L g4851 ( 
.A1(n_4757),
.A2(n_592),
.B(n_593),
.Y(n_4851)
);

OAI22xp5_ASAP7_75t_SL g4852 ( 
.A1(n_4794),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4750),
.B(n_594),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4796),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4761),
.Y(n_4855)
);

NAND2xp33_ASAP7_75t_L g4856 ( 
.A(n_4768),
.B(n_595),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4845),
.Y(n_4857)
);

INVx1_ASAP7_75t_SL g4858 ( 
.A(n_4850),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4845),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4840),
.Y(n_4860)
);

NOR2xp33_ASAP7_75t_L g4861 ( 
.A(n_4842),
.B(n_599),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4808),
.Y(n_4862)
);

OAI21xp33_ASAP7_75t_L g4863 ( 
.A1(n_4803),
.A2(n_609),
.B(n_599),
.Y(n_4863)
);

NAND2x1_ASAP7_75t_L g4864 ( 
.A(n_4800),
.B(n_601),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4809),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4821),
.B(n_601),
.Y(n_4866)
);

OR2x2_ASAP7_75t_L g4867 ( 
.A(n_4854),
.B(n_602),
.Y(n_4867)
);

AOI32xp33_ASAP7_75t_L g4868 ( 
.A1(n_4851),
.A2(n_604),
.A3(n_602),
.B1(n_603),
.B2(n_605),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4843),
.Y(n_4869)
);

NOR2xp33_ASAP7_75t_L g4870 ( 
.A(n_4811),
.B(n_604),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4853),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4852),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4817),
.Y(n_4873)
);

XOR2x2_ASAP7_75t_L g4874 ( 
.A(n_4839),
.B(n_4814),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4820),
.B(n_605),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4856),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4816),
.B(n_606),
.Y(n_4877)
);

OAI21xp5_ASAP7_75t_SL g4878 ( 
.A1(n_4806),
.A2(n_606),
.B(n_608),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4801),
.B(n_608),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4812),
.Y(n_4880)
);

OAI31xp33_ASAP7_75t_L g4881 ( 
.A1(n_4804),
.A2(n_612),
.A3(n_610),
.B(n_611),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_SL g4882 ( 
.A(n_4810),
.B(n_610),
.Y(n_4882)
);

NAND2xp33_ASAP7_75t_L g4883 ( 
.A(n_4832),
.B(n_611),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4819),
.Y(n_4884)
);

NOR2x1_ASAP7_75t_L g4885 ( 
.A(n_4838),
.B(n_612),
.Y(n_4885)
);

AOI22xp5_ASAP7_75t_L g4886 ( 
.A1(n_4807),
.A2(n_616),
.B1(n_613),
.B2(n_615),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4841),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4802),
.B(n_613),
.Y(n_4888)
);

AOI221xp5_ASAP7_75t_L g4889 ( 
.A1(n_4799),
.A2(n_4847),
.B1(n_4855),
.B2(n_4848),
.C(n_4844),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4829),
.Y(n_4890)
);

AND2x4_ASAP7_75t_SL g4891 ( 
.A(n_4831),
.B(n_615),
.Y(n_4891)
);

INVx1_ASAP7_75t_SL g4892 ( 
.A(n_4849),
.Y(n_4892)
);

XOR2x2_ASAP7_75t_L g4893 ( 
.A(n_4815),
.B(n_616),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4834),
.B(n_617),
.Y(n_4894)
);

A2O1A1Ixp33_ASAP7_75t_SL g4895 ( 
.A1(n_4823),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4837),
.B(n_618),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4826),
.B(n_619),
.Y(n_4897)
);

NOR2x1_ASAP7_75t_L g4898 ( 
.A(n_4824),
.B(n_620),
.Y(n_4898)
);

AOI22xp5_ASAP7_75t_L g4899 ( 
.A1(n_4822),
.A2(n_4828),
.B1(n_4813),
.B2(n_4798),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4818),
.B(n_620),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4827),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4835),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4846),
.B(n_621),
.Y(n_4903)
);

INVx1_ASAP7_75t_SL g4904 ( 
.A(n_4825),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4805),
.Y(n_4905)
);

AOI221x1_ASAP7_75t_L g4906 ( 
.A1(n_4833),
.A2(n_623),
.B1(n_626),
.B2(n_622),
.C(n_625),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4836),
.B(n_621),
.Y(n_4907)
);

XNOR2xp5_ASAP7_75t_L g4908 ( 
.A(n_4830),
.B(n_625),
.Y(n_4908)
);

OAI222xp33_ASAP7_75t_L g4909 ( 
.A1(n_4842),
.A2(n_627),
.B1(n_629),
.B2(n_622),
.C1(n_626),
.C2(n_628),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4800),
.B(n_627),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4845),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4845),
.B(n_629),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4800),
.B(n_630),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4845),
.B(n_630),
.Y(n_4914)
);

AOI21xp5_ASAP7_75t_L g4915 ( 
.A1(n_4803),
.A2(n_632),
.B(n_633),
.Y(n_4915)
);

AOI22xp5_ASAP7_75t_L g4916 ( 
.A1(n_4803),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_4916)
);

AND2x4_ASAP7_75t_L g4917 ( 
.A(n_4845),
.B(n_635),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4845),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4800),
.B(n_636),
.Y(n_4919)
);

AND3x1_ASAP7_75t_L g4920 ( 
.A(n_4803),
.B(n_637),
.C(n_638),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4845),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4803),
.A2(n_639),
.B(n_640),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4845),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4845),
.B(n_639),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4845),
.B(n_642),
.Y(n_4925)
);

AOI211xp5_ASAP7_75t_SL g4926 ( 
.A1(n_4803),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_4926)
);

O2A1O1Ixp33_ASAP7_75t_L g4927 ( 
.A1(n_4803),
.A2(n_654),
.B(n_665),
.C(n_644),
.Y(n_4927)
);

OR2x2_ASAP7_75t_L g4928 ( 
.A(n_4845),
.B(n_646),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4845),
.B(n_646),
.Y(n_4929)
);

AOI22xp33_ASAP7_75t_SL g4930 ( 
.A1(n_4839),
.A2(n_650),
.B1(n_647),
.B2(n_648),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4845),
.B(n_650),
.Y(n_4931)
);

NAND5xp2_ASAP7_75t_L g4932 ( 
.A(n_4815),
.B(n_653),
.C(n_651),
.D(n_652),
.E(n_656),
.Y(n_4932)
);

OAI211xp5_ASAP7_75t_SL g4933 ( 
.A1(n_4803),
.A2(n_656),
.B(n_652),
.C(n_653),
.Y(n_4933)
);

AOI211x1_ASAP7_75t_L g4934 ( 
.A1(n_4803),
.A2(n_661),
.B(n_657),
.C(n_660),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4845),
.Y(n_4935)
);

NOR2x1_ASAP7_75t_L g4936 ( 
.A(n_4814),
.B(n_660),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4800),
.B(n_662),
.Y(n_4937)
);

INVxp67_ASAP7_75t_L g4938 ( 
.A(n_4807),
.Y(n_4938)
);

INVx1_ASAP7_75t_SL g4939 ( 
.A(n_4850),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4845),
.B(n_662),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4845),
.B(n_663),
.Y(n_4941)
);

INVx1_ASAP7_75t_SL g4942 ( 
.A(n_4850),
.Y(n_4942)
);

OAI22xp5_ASAP7_75t_L g4943 ( 
.A1(n_4839),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4845),
.B(n_666),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4845),
.B(n_667),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_4845),
.B(n_668),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4845),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4845),
.Y(n_4948)
);

INVx1_ASAP7_75t_SL g4949 ( 
.A(n_4891),
.Y(n_4949)
);

NAND2xp33_ASAP7_75t_SL g4950 ( 
.A(n_4864),
.B(n_669),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4928),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4859),
.Y(n_4952)
);

NOR3xp33_ASAP7_75t_L g4953 ( 
.A(n_4938),
.B(n_669),
.C(n_670),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4857),
.B(n_4947),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4911),
.B(n_672),
.Y(n_4955)
);

O2A1O1Ixp5_ASAP7_75t_SL g4956 ( 
.A1(n_4918),
.A2(n_675),
.B(n_673),
.C(n_674),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4921),
.B(n_673),
.Y(n_4957)
);

NAND3xp33_ASAP7_75t_L g4958 ( 
.A(n_4926),
.B(n_674),
.C(n_677),
.Y(n_4958)
);

AOI21xp33_ASAP7_75t_L g4959 ( 
.A1(n_4883),
.A2(n_677),
.B(n_678),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_4923),
.B(n_679),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4935),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4948),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4887),
.B(n_679),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4858),
.B(n_680),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4917),
.Y(n_4965)
);

NOR2xp33_ASAP7_75t_L g4966 ( 
.A(n_4932),
.B(n_680),
.Y(n_4966)
);

XOR2xp5_ASAP7_75t_L g4967 ( 
.A(n_4874),
.B(n_681),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4917),
.Y(n_4968)
);

NOR2xp33_ASAP7_75t_L g4969 ( 
.A(n_4939),
.B(n_681),
.Y(n_4969)
);

OR2x2_ASAP7_75t_L g4970 ( 
.A(n_4942),
.B(n_4880),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4890),
.B(n_4872),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4912),
.Y(n_4972)
);

INVx3_ASAP7_75t_L g4973 ( 
.A(n_4873),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4914),
.Y(n_4974)
);

AND2x4_ASAP7_75t_L g4975 ( 
.A(n_4898),
.B(n_4860),
.Y(n_4975)
);

INVxp67_ASAP7_75t_L g4976 ( 
.A(n_4885),
.Y(n_4976)
);

OR2x2_ASAP7_75t_L g4977 ( 
.A(n_4892),
.B(n_682),
.Y(n_4977)
);

INVxp33_ASAP7_75t_SL g4978 ( 
.A(n_4899),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4930),
.B(n_4934),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4924),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_4893),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4925),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4867),
.Y(n_4983)
);

OAI21xp5_ASAP7_75t_SL g4984 ( 
.A1(n_4916),
.A2(n_4868),
.B(n_4878),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4875),
.Y(n_4985)
);

OAI211xp5_ASAP7_75t_L g4986 ( 
.A1(n_4863),
.A2(n_693),
.B(n_702),
.C(n_682),
.Y(n_4986)
);

NOR2xp33_ASAP7_75t_L g4987 ( 
.A(n_4933),
.B(n_684),
.Y(n_4987)
);

CKINVDCx20_ASAP7_75t_R g4988 ( 
.A(n_4905),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4929),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4931),
.Y(n_4990)
);

BUFx4f_ASAP7_75t_SL g4991 ( 
.A(n_4904),
.Y(n_4991)
);

OR2x2_ASAP7_75t_L g4992 ( 
.A(n_4866),
.B(n_684),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4886),
.B(n_685),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4876),
.B(n_685),
.Y(n_4994)
);

AOI21xp33_ASAP7_75t_L g4995 ( 
.A1(n_4927),
.A2(n_687),
.B(n_688),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4940),
.Y(n_4996)
);

OAI22xp33_ASAP7_75t_SL g4997 ( 
.A1(n_4882),
.A2(n_692),
.B1(n_689),
.B2(n_690),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4941),
.Y(n_4998)
);

AND2x2_ASAP7_75t_L g4999 ( 
.A(n_4910),
.B(n_690),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4944),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4913),
.B(n_692),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4919),
.B(n_4937),
.Y(n_5002)
);

HB1xp67_ASAP7_75t_L g5003 ( 
.A(n_4936),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4884),
.B(n_694),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4945),
.Y(n_5005)
);

OR2x2_ASAP7_75t_L g5006 ( 
.A(n_4877),
.B(n_4943),
.Y(n_5006)
);

INVx2_ASAP7_75t_L g5007 ( 
.A(n_4894),
.Y(n_5007)
);

INVxp67_ASAP7_75t_L g5008 ( 
.A(n_4870),
.Y(n_5008)
);

AND2x2_ASAP7_75t_SL g5009 ( 
.A(n_4920),
.B(n_695),
.Y(n_5009)
);

NOR2xp33_ASAP7_75t_L g5010 ( 
.A(n_4879),
.B(n_696),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4946),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4908),
.Y(n_5012)
);

OR2x2_ASAP7_75t_L g5013 ( 
.A(n_4896),
.B(n_696),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4900),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4915),
.B(n_697),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4903),
.Y(n_5016)
);

INVx3_ASAP7_75t_L g5017 ( 
.A(n_4862),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4922),
.B(n_697),
.Y(n_5018)
);

AOI21xp5_ASAP7_75t_L g5019 ( 
.A1(n_4895),
.A2(n_698),
.B(n_699),
.Y(n_5019)
);

INVx2_ASAP7_75t_SL g5020 ( 
.A(n_4865),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4888),
.Y(n_5021)
);

AND2x2_ASAP7_75t_L g5022 ( 
.A(n_4869),
.B(n_699),
.Y(n_5022)
);

AOI22xp33_ASAP7_75t_R g5023 ( 
.A1(n_4871),
.A2(n_703),
.B1(n_700),
.B2(n_702),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4897),
.Y(n_5024)
);

OAI21xp33_ASAP7_75t_L g5025 ( 
.A1(n_4889),
.A2(n_4861),
.B(n_4902),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4881),
.B(n_700),
.Y(n_5026)
);

OAI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4907),
.A2(n_703),
.B(n_704),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4906),
.B(n_704),
.Y(n_5028)
);

AOI21xp33_ASAP7_75t_SL g5029 ( 
.A1(n_4901),
.A2(n_4909),
.B(n_705),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4928),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4928),
.Y(n_5031)
);

INVx2_ASAP7_75t_SL g5032 ( 
.A(n_4891),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4928),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_4859),
.B(n_706),
.Y(n_5034)
);

AOI22xp33_ASAP7_75t_SL g5035 ( 
.A1(n_4860),
.A2(n_709),
.B1(n_707),
.B2(n_708),
.Y(n_5035)
);

INVx1_ASAP7_75t_SL g5036 ( 
.A(n_4891),
.Y(n_5036)
);

NOR3x1_ASAP7_75t_L g5037 ( 
.A(n_4958),
.B(n_707),
.C(n_709),
.Y(n_5037)
);

AOI31xp33_ASAP7_75t_L g5038 ( 
.A1(n_4976),
.A2(n_718),
.A3(n_727),
.B(n_710),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4965),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_5009),
.B(n_710),
.Y(n_5040)
);

OA22x2_ASAP7_75t_L g5041 ( 
.A1(n_4967),
.A2(n_713),
.B1(n_711),
.B2(n_712),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4968),
.B(n_711),
.Y(n_5042)
);

AOI221xp5_ASAP7_75t_L g5043 ( 
.A1(n_5029),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.C(n_716),
.Y(n_5043)
);

AOI21xp5_ASAP7_75t_L g5044 ( 
.A1(n_4950),
.A2(n_716),
.B(n_717),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4977),
.Y(n_5045)
);

OAI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_5019),
.A2(n_719),
.B(n_718),
.Y(n_5046)
);

AOI22xp5_ASAP7_75t_L g5047 ( 
.A1(n_4988),
.A2(n_721),
.B1(n_717),
.B2(n_720),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_5032),
.B(n_720),
.Y(n_5048)
);

NOR2x1p5_ASAP7_75t_L g5049 ( 
.A(n_4973),
.B(n_722),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4949),
.B(n_723),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_5036),
.B(n_723),
.Y(n_5051)
);

INVx1_ASAP7_75t_SL g5052 ( 
.A(n_4991),
.Y(n_5052)
);

NOR3xp33_ASAP7_75t_L g5053 ( 
.A(n_5025),
.B(n_727),
.C(n_725),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4999),
.Y(n_5054)
);

AOI211x1_ASAP7_75t_L g5055 ( 
.A1(n_4995),
.A2(n_4959),
.B(n_4971),
.C(n_4979),
.Y(n_5055)
);

NOR3xp33_ASAP7_75t_L g5056 ( 
.A(n_4970),
.B(n_728),
.C(n_725),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4966),
.B(n_5035),
.Y(n_5057)
);

OAI22xp5_ASAP7_75t_L g5058 ( 
.A1(n_4978),
.A2(n_729),
.B1(n_724),
.B2(n_728),
.Y(n_5058)
);

NOR2xp67_ASAP7_75t_L g5059 ( 
.A(n_5003),
.B(n_729),
.Y(n_5059)
);

OAI31xp33_ASAP7_75t_L g5060 ( 
.A1(n_4997),
.A2(n_731),
.A3(n_724),
.B(n_730),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_5004),
.Y(n_5061)
);

OAI211xp5_ASAP7_75t_L g5062 ( 
.A1(n_4984),
.A2(n_732),
.B(n_730),
.C(n_731),
.Y(n_5062)
);

NOR3xp33_ASAP7_75t_L g5063 ( 
.A(n_5002),
.B(n_735),
.C(n_734),
.Y(n_5063)
);

AOI22xp5_ASAP7_75t_L g5064 ( 
.A1(n_4981),
.A2(n_737),
.B1(n_732),
.B2(n_736),
.Y(n_5064)
);

AOI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4987),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4975),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4975),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4985),
.B(n_738),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4952),
.B(n_739),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4969),
.B(n_740),
.Y(n_5070)
);

OA211x2_ASAP7_75t_L g5071 ( 
.A1(n_5028),
.A2(n_742),
.B(n_740),
.C(n_741),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_5007),
.B(n_5022),
.Y(n_5072)
);

NOR3xp33_ASAP7_75t_L g5073 ( 
.A(n_5026),
.B(n_4963),
.C(n_4954),
.Y(n_5073)
);

NOR3xp33_ASAP7_75t_L g5074 ( 
.A(n_5012),
.B(n_743),
.C(n_742),
.Y(n_5074)
);

AOI211xp5_ASAP7_75t_L g5075 ( 
.A1(n_4986),
.A2(n_744),
.B(n_741),
.C(n_743),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4964),
.Y(n_5076)
);

OAI21xp33_ASAP7_75t_SL g5077 ( 
.A1(n_5020),
.A2(n_744),
.B(n_745),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_5001),
.Y(n_5078)
);

AOI211xp5_ASAP7_75t_L g5079 ( 
.A1(n_4961),
.A2(n_747),
.B(n_745),
.C(n_746),
.Y(n_5079)
);

AOI211xp5_ASAP7_75t_L g5080 ( 
.A1(n_4962),
.A2(n_748),
.B(n_746),
.C(n_747),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_4983),
.B(n_5014),
.Y(n_5081)
);

AOI211xp5_ASAP7_75t_L g5082 ( 
.A1(n_5027),
.A2(n_750),
.B(n_748),
.C(n_749),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4953),
.B(n_749),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_4951),
.B(n_751),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_SL g5085 ( 
.A(n_5017),
.B(n_751),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4994),
.Y(n_5086)
);

NOR3x1_ASAP7_75t_L g5087 ( 
.A(n_5015),
.B(n_752),
.C(n_753),
.Y(n_5087)
);

NAND2xp33_ASAP7_75t_SL g5088 ( 
.A(n_5030),
.B(n_753),
.Y(n_5088)
);

AO21x1_ASAP7_75t_L g5089 ( 
.A1(n_4955),
.A2(n_754),
.B(n_755),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4992),
.Y(n_5090)
);

NOR2x1_ASAP7_75t_L g5091 ( 
.A(n_5031),
.B(n_756),
.Y(n_5091)
);

NOR2x1_ASAP7_75t_L g5092 ( 
.A(n_5033),
.B(n_756),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_5010),
.B(n_757),
.Y(n_5093)
);

NOR3xp33_ASAP7_75t_L g5094 ( 
.A(n_5008),
.B(n_759),
.C(n_758),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_5034),
.Y(n_5095)
);

OA22x2_ASAP7_75t_L g5096 ( 
.A1(n_4957),
.A2(n_760),
.B1(n_757),
.B2(n_758),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4960),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_SL g5098 ( 
.A(n_5018),
.B(n_760),
.Y(n_5098)
);

AOI21xp5_ASAP7_75t_L g5099 ( 
.A1(n_4993),
.A2(n_5006),
.B(n_5013),
.Y(n_5099)
);

OAI21xp33_ASAP7_75t_L g5100 ( 
.A1(n_5016),
.A2(n_761),
.B(n_762),
.Y(n_5100)
);

AO22x2_ASAP7_75t_L g5101 ( 
.A1(n_5024),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_5101)
);

XNOR2xp5_ASAP7_75t_L g5102 ( 
.A(n_5023),
.B(n_763),
.Y(n_5102)
);

NOR2x1_ASAP7_75t_L g5103 ( 
.A(n_4972),
.B(n_765),
.Y(n_5103)
);

NOR3x1_ASAP7_75t_L g5104 ( 
.A(n_4974),
.B(n_4982),
.C(n_4980),
.Y(n_5104)
);

NOR3xp33_ASAP7_75t_L g5105 ( 
.A(n_4989),
.B(n_767),
.C(n_766),
.Y(n_5105)
);

AOI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_4990),
.A2(n_767),
.B1(n_765),
.B2(n_766),
.Y(n_5106)
);

AOI21xp5_ASAP7_75t_L g5107 ( 
.A1(n_4996),
.A2(n_768),
.B(n_769),
.Y(n_5107)
);

INVx3_ASAP7_75t_L g5108 ( 
.A(n_4998),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_5000),
.A2(n_5011),
.B(n_5005),
.Y(n_5109)
);

AOI211x1_ASAP7_75t_L g5110 ( 
.A1(n_5021),
.A2(n_771),
.B(n_768),
.C(n_770),
.Y(n_5110)
);

AOI21xp5_ASAP7_75t_L g5111 ( 
.A1(n_4956),
.A2(n_770),
.B(n_772),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_5009),
.B(n_772),
.Y(n_5112)
);

AOI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_4950),
.A2(n_773),
.B(n_774),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_SL g5114 ( 
.A1(n_4975),
.A2(n_774),
.B(n_775),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4965),
.Y(n_5115)
);

NOR2xp33_ASAP7_75t_SL g5116 ( 
.A(n_5009),
.B(n_776),
.Y(n_5116)
);

AOI211x1_ASAP7_75t_L g5117 ( 
.A1(n_4995),
.A2(n_779),
.B(n_777),
.C(n_778),
.Y(n_5117)
);

NAND2xp5_ASAP7_75t_L g5118 ( 
.A(n_5009),
.B(n_778),
.Y(n_5118)
);

NOR2x1_ASAP7_75t_L g5119 ( 
.A(n_5028),
.B(n_779),
.Y(n_5119)
);

O2A1O1Ixp33_ASAP7_75t_SL g5120 ( 
.A1(n_4976),
.A2(n_789),
.B(n_798),
.C(n_780),
.Y(n_5120)
);

AOI22xp5_ASAP7_75t_L g5121 ( 
.A1(n_4988),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_5121)
);

NOR3xp33_ASAP7_75t_L g5122 ( 
.A(n_5025),
.B(n_785),
.C(n_784),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4965),
.Y(n_5123)
);

INVx1_ASAP7_75t_SL g5124 ( 
.A(n_5088),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_5041),
.Y(n_5125)
);

XOR2x2_ASAP7_75t_L g5126 ( 
.A(n_5052),
.B(n_783),
.Y(n_5126)
);

XNOR2x1_ASAP7_75t_L g5127 ( 
.A(n_5071),
.B(n_784),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5091),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_SL g5129 ( 
.A(n_5116),
.B(n_785),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_5092),
.Y(n_5130)
);

NOR2x1_ASAP7_75t_L g5131 ( 
.A(n_5114),
.B(n_787),
.Y(n_5131)
);

XOR2x2_ASAP7_75t_L g5132 ( 
.A(n_5119),
.B(n_787),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5089),
.Y(n_5133)
);

CKINVDCx16_ASAP7_75t_R g5134 ( 
.A(n_5081),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5096),
.Y(n_5135)
);

OAI21xp33_ASAP7_75t_L g5136 ( 
.A1(n_5057),
.A2(n_788),
.B(n_790),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_5059),
.Y(n_5137)
);

NOR2x1_ASAP7_75t_L g5138 ( 
.A(n_5103),
.B(n_788),
.Y(n_5138)
);

A2O1A1Ixp33_ASAP7_75t_L g5139 ( 
.A1(n_5044),
.A2(n_793),
.B(n_790),
.C(n_791),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5040),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5112),
.Y(n_5141)
);

AND2x2_ASAP7_75t_L g5142 ( 
.A(n_5039),
.B(n_5115),
.Y(n_5142)
);

AOI22xp5_ASAP7_75t_L g5143 ( 
.A1(n_5123),
.A2(n_5073),
.B1(n_5122),
.B2(n_5053),
.Y(n_5143)
);

INVx2_ASAP7_75t_SL g5144 ( 
.A(n_5049),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5118),
.Y(n_5145)
);

NAND3x2_ASAP7_75t_L g5146 ( 
.A(n_5066),
.B(n_791),
.C(n_794),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_5120),
.Y(n_5147)
);

AOI322xp5_ASAP7_75t_L g5148 ( 
.A1(n_5067),
.A2(n_800),
.A3(n_799),
.B1(n_796),
.B2(n_794),
.C1(n_795),
.C2(n_797),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_5101),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_5113),
.B(n_797),
.Y(n_5150)
);

XNOR2x1_ASAP7_75t_L g5151 ( 
.A(n_5102),
.B(n_799),
.Y(n_5151)
);

INVx1_ASAP7_75t_SL g5152 ( 
.A(n_5084),
.Y(n_5152)
);

AOI22xp5_ASAP7_75t_L g5153 ( 
.A1(n_5054),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_5101),
.Y(n_5154)
);

INVx1_ASAP7_75t_SL g5155 ( 
.A(n_5068),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_5111),
.B(n_802),
.Y(n_5156)
);

NOR2x1_ASAP7_75t_L g5157 ( 
.A(n_5038),
.B(n_803),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_5046),
.B(n_805),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5050),
.Y(n_5159)
);

OAI21xp5_ASAP7_75t_L g5160 ( 
.A1(n_5077),
.A2(n_805),
.B(n_806),
.Y(n_5160)
);

AOI32xp33_ASAP7_75t_L g5161 ( 
.A1(n_5043),
.A2(n_809),
.A3(n_811),
.B1(n_808),
.B2(n_810),
.Y(n_5161)
);

INVx2_ASAP7_75t_SL g5162 ( 
.A(n_5108),
.Y(n_5162)
);

XNOR2x1_ASAP7_75t_L g5163 ( 
.A(n_5065),
.B(n_806),
.Y(n_5163)
);

BUFx3_ASAP7_75t_L g5164 ( 
.A(n_5061),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5110),
.B(n_809),
.Y(n_5165)
);

OAI22xp33_ASAP7_75t_SL g5166 ( 
.A1(n_5051),
.A2(n_814),
.B1(n_811),
.B2(n_812),
.Y(n_5166)
);

NOR2x1_ASAP7_75t_L g5167 ( 
.A(n_5062),
.B(n_814),
.Y(n_5167)
);

NOR3xp33_ASAP7_75t_L g5168 ( 
.A(n_5072),
.B(n_815),
.C(n_816),
.Y(n_5168)
);

OAI21xp5_ASAP7_75t_L g5169 ( 
.A1(n_5109),
.A2(n_5048),
.B(n_5099),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5079),
.B(n_815),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5080),
.B(n_816),
.Y(n_5171)
);

INVx2_ASAP7_75t_L g5172 ( 
.A(n_5087),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5060),
.B(n_817),
.Y(n_5173)
);

HB1xp67_ASAP7_75t_L g5174 ( 
.A(n_5058),
.Y(n_5174)
);

AOI22xp33_ASAP7_75t_L g5175 ( 
.A1(n_5045),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_5175)
);

OAI21xp5_ASAP7_75t_L g5176 ( 
.A1(n_5042),
.A2(n_818),
.B(n_820),
.Y(n_5176)
);

AND2x2_ASAP7_75t_L g5177 ( 
.A(n_5037),
.B(n_820),
.Y(n_5177)
);

AOI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_5056),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_5178)
);

AOI221xp5_ASAP7_75t_L g5179 ( 
.A1(n_5055),
.A2(n_824),
.B1(n_821),
.B2(n_823),
.C(n_825),
.Y(n_5179)
);

XOR2xp5_ASAP7_75t_L g5180 ( 
.A(n_5064),
.B(n_824),
.Y(n_5180)
);

AOI211x1_ASAP7_75t_SL g5181 ( 
.A1(n_5098),
.A2(n_828),
.B(n_825),
.C(n_827),
.Y(n_5181)
);

NOR3xp33_ASAP7_75t_L g5182 ( 
.A(n_5108),
.B(n_828),
.C(n_829),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5069),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_5070),
.Y(n_5184)
);

NOR2xp33_ASAP7_75t_L g5185 ( 
.A(n_5100),
.B(n_829),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5083),
.Y(n_5186)
);

NOR3xp33_ASAP7_75t_L g5187 ( 
.A(n_5090),
.B(n_830),
.C(n_831),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_5107),
.B(n_831),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5085),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_5093),
.Y(n_5190)
);

NAND3xp33_ASAP7_75t_L g5191 ( 
.A(n_5075),
.B(n_832),
.C(n_833),
.Y(n_5191)
);

OAI22xp33_ASAP7_75t_L g5192 ( 
.A1(n_5121),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.Y(n_5192)
);

AOI21xp33_ASAP7_75t_L g5193 ( 
.A1(n_5076),
.A2(n_834),
.B(n_836),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_SL g5194 ( 
.A(n_5063),
.B(n_836),
.Y(n_5194)
);

INVx1_ASAP7_75t_SL g5195 ( 
.A(n_5047),
.Y(n_5195)
);

O2A1O1Ixp5_ASAP7_75t_SL g5196 ( 
.A1(n_5086),
.A2(n_842),
.B(n_840),
.C(n_841),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5117),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5105),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5094),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5074),
.Y(n_5200)
);

AND2x2_ASAP7_75t_L g5201 ( 
.A(n_5134),
.B(n_5104),
.Y(n_5201)
);

OAI22xp5_ASAP7_75t_SL g5202 ( 
.A1(n_5147),
.A2(n_5082),
.B1(n_5078),
.B2(n_5095),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5131),
.Y(n_5203)
);

AOI22xp5_ASAP7_75t_L g5204 ( 
.A1(n_5125),
.A2(n_5097),
.B1(n_5106),
.B2(n_844),
.Y(n_5204)
);

NOR4xp25_ASAP7_75t_L g5205 ( 
.A(n_5124),
.B(n_844),
.C(n_841),
.D(n_843),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5127),
.Y(n_5206)
);

NOR2x1_ASAP7_75t_L g5207 ( 
.A(n_5138),
.B(n_845),
.Y(n_5207)
);

AO22x2_ASAP7_75t_SL g5208 ( 
.A1(n_5133),
.A2(n_847),
.B1(n_845),
.B2(n_846),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_5149),
.B(n_846),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_5126),
.Y(n_5210)
);

NOR2x1_ASAP7_75t_L g5211 ( 
.A(n_5128),
.B(n_847),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_5154),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5157),
.Y(n_5213)
);

NOR2x1_ASAP7_75t_L g5214 ( 
.A(n_5130),
.B(n_848),
.Y(n_5214)
);

NOR2x1_ASAP7_75t_L g5215 ( 
.A(n_5137),
.B(n_848),
.Y(n_5215)
);

AO22x2_ASAP7_75t_L g5216 ( 
.A1(n_5162),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5177),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5142),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_5132),
.Y(n_5219)
);

XNOR2x1_ASAP7_75t_L g5220 ( 
.A(n_5151),
.B(n_850),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5156),
.Y(n_5221)
);

AOI22xp5_ASAP7_75t_L g5222 ( 
.A1(n_5135),
.A2(n_853),
.B1(n_851),
.B2(n_852),
.Y(n_5222)
);

AOI22xp5_ASAP7_75t_L g5223 ( 
.A1(n_5152),
.A2(n_857),
.B1(n_854),
.B2(n_856),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5165),
.Y(n_5224)
);

HB1xp67_ASAP7_75t_L g5225 ( 
.A(n_5160),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5150),
.Y(n_5226)
);

AO22x2_ASAP7_75t_L g5227 ( 
.A1(n_5144),
.A2(n_858),
.B1(n_854),
.B2(n_856),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5167),
.Y(n_5228)
);

AOI31xp33_ASAP7_75t_L g5229 ( 
.A1(n_5129),
.A2(n_866),
.A3(n_874),
.B(n_858),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5174),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5182),
.B(n_859),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_5173),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5188),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_5187),
.B(n_859),
.Y(n_5234)
);

OA22x2_ASAP7_75t_L g5235 ( 
.A1(n_5143),
.A2(n_862),
.B1(n_860),
.B2(n_861),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5164),
.Y(n_5236)
);

AOI22xp5_ASAP7_75t_L g5237 ( 
.A1(n_5197),
.A2(n_5195),
.B1(n_5155),
.B2(n_5172),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_SL g5238 ( 
.A(n_5166),
.B(n_860),
.Y(n_5238)
);

OA22x2_ASAP7_75t_L g5239 ( 
.A1(n_5180),
.A2(n_865),
.B1(n_863),
.B2(n_864),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5170),
.Y(n_5240)
);

OA22x2_ASAP7_75t_L g5241 ( 
.A1(n_5178),
.A2(n_868),
.B1(n_864),
.B2(n_867),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_SL g5242 ( 
.A(n_5179),
.B(n_867),
.Y(n_5242)
);

AOI31xp33_ASAP7_75t_L g5243 ( 
.A1(n_5169),
.A2(n_871),
.A3(n_869),
.B(n_870),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_SL g5244 ( 
.A(n_5192),
.B(n_869),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_5139),
.B(n_870),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_5171),
.Y(n_5246)
);

HB1xp67_ASAP7_75t_L g5247 ( 
.A(n_5181),
.Y(n_5247)
);

OAI22xp5_ASAP7_75t_SL g5248 ( 
.A1(n_5191),
.A2(n_874),
.B1(n_872),
.B2(n_873),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5158),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5136),
.Y(n_5250)
);

AO22x1_ASAP7_75t_L g5251 ( 
.A1(n_5168),
.A2(n_877),
.B1(n_875),
.B2(n_876),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5185),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_5163),
.Y(n_5253)
);

OA22x2_ASAP7_75t_L g5254 ( 
.A1(n_5189),
.A2(n_878),
.B1(n_876),
.B2(n_877),
.Y(n_5254)
);

AOI22xp5_ASAP7_75t_L g5255 ( 
.A1(n_5200),
.A2(n_882),
.B1(n_878),
.B2(n_881),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_5176),
.Y(n_5256)
);

OAI22xp33_ASAP7_75t_L g5257 ( 
.A1(n_5243),
.A2(n_5198),
.B1(n_5199),
.B2(n_5159),
.Y(n_5257)
);

OAI221xp5_ASAP7_75t_L g5258 ( 
.A1(n_5237),
.A2(n_5161),
.B1(n_5205),
.B2(n_5206),
.C(n_5212),
.Y(n_5258)
);

NOR2xp33_ASAP7_75t_R g5259 ( 
.A(n_5203),
.B(n_5140),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_5208),
.Y(n_5260)
);

OAI211xp5_ASAP7_75t_SL g5261 ( 
.A1(n_5230),
.A2(n_5145),
.B(n_5141),
.C(n_5186),
.Y(n_5261)
);

NOR3xp33_ASAP7_75t_L g5262 ( 
.A(n_5202),
.B(n_5183),
.C(n_5184),
.Y(n_5262)
);

AOI322xp5_ASAP7_75t_L g5263 ( 
.A1(n_5201),
.A2(n_5194),
.A3(n_5190),
.B1(n_5193),
.B2(n_5175),
.C1(n_5153),
.C2(n_5146),
.Y(n_5263)
);

NAND3xp33_ASAP7_75t_L g5264 ( 
.A(n_5207),
.B(n_5196),
.C(n_5148),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5254),
.Y(n_5265)
);

AOI211xp5_ASAP7_75t_L g5266 ( 
.A1(n_5248),
.A2(n_5251),
.B(n_5236),
.C(n_5218),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_5215),
.B(n_882),
.Y(n_5267)
);

XNOR2xp5_ASAP7_75t_L g5268 ( 
.A(n_5220),
.B(n_883),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_5222),
.B(n_5211),
.Y(n_5269)
);

HB1xp67_ASAP7_75t_L g5270 ( 
.A(n_5216),
.Y(n_5270)
);

OR2x2_ASAP7_75t_L g5271 ( 
.A(n_5209),
.B(n_5213),
.Y(n_5271)
);

AOI221xp5_ASAP7_75t_L g5272 ( 
.A1(n_5228),
.A2(n_885),
.B1(n_883),
.B2(n_884),
.C(n_886),
.Y(n_5272)
);

NAND2xp33_ASAP7_75t_SL g5273 ( 
.A(n_5247),
.B(n_885),
.Y(n_5273)
);

OAI211xp5_ASAP7_75t_SL g5274 ( 
.A1(n_5204),
.A2(n_888),
.B(n_886),
.C(n_887),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_5235),
.Y(n_5275)
);

NOR2xp33_ASAP7_75t_L g5276 ( 
.A(n_5229),
.B(n_887),
.Y(n_5276)
);

INVx1_ASAP7_75t_SL g5277 ( 
.A(n_5214),
.Y(n_5277)
);

NAND3xp33_ASAP7_75t_L g5278 ( 
.A(n_5238),
.B(n_889),
.C(n_890),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_5217),
.B(n_889),
.Y(n_5279)
);

OAI211xp5_ASAP7_75t_SL g5280 ( 
.A1(n_5242),
.A2(n_892),
.B(n_890),
.C(n_891),
.Y(n_5280)
);

NAND2xp5_ASAP7_75t_SL g5281 ( 
.A(n_5239),
.B(n_891),
.Y(n_5281)
);

OAI21xp5_ASAP7_75t_SL g5282 ( 
.A1(n_5210),
.A2(n_892),
.B(n_894),
.Y(n_5282)
);

AOI22xp5_ASAP7_75t_L g5283 ( 
.A1(n_5219),
.A2(n_897),
.B1(n_895),
.B2(n_896),
.Y(n_5283)
);

CKINVDCx20_ASAP7_75t_R g5284 ( 
.A(n_5225),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5241),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_5223),
.B(n_895),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_5255),
.B(n_896),
.Y(n_5287)
);

AOI22xp33_ASAP7_75t_L g5288 ( 
.A1(n_5224),
.A2(n_899),
.B1(n_897),
.B2(n_898),
.Y(n_5288)
);

NAND3xp33_ASAP7_75t_L g5289 ( 
.A(n_5231),
.B(n_898),
.C(n_899),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5216),
.Y(n_5290)
);

NAND2xp33_ASAP7_75t_SL g5291 ( 
.A(n_5245),
.B(n_900),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5270),
.Y(n_5292)
);

INVxp67_ASAP7_75t_L g5293 ( 
.A(n_5276),
.Y(n_5293)
);

OAI211xp5_ASAP7_75t_SL g5294 ( 
.A1(n_5263),
.A2(n_5250),
.B(n_5253),
.C(n_5256),
.Y(n_5294)
);

NOR2xp67_ASAP7_75t_L g5295 ( 
.A(n_5290),
.B(n_5234),
.Y(n_5295)
);

AND2x4_ASAP7_75t_L g5296 ( 
.A(n_5262),
.B(n_5249),
.Y(n_5296)
);

XOR2xp5_ASAP7_75t_L g5297 ( 
.A(n_5268),
.B(n_5284),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_5279),
.Y(n_5298)
);

BUFx4f_ASAP7_75t_L g5299 ( 
.A(n_5271),
.Y(n_5299)
);

NOR3xp33_ASAP7_75t_L g5300 ( 
.A(n_5261),
.B(n_5221),
.C(n_5232),
.Y(n_5300)
);

NAND2xp33_ASAP7_75t_L g5301 ( 
.A(n_5277),
.B(n_5260),
.Y(n_5301)
);

NAND4xp75_ASAP7_75t_L g5302 ( 
.A(n_5285),
.B(n_5252),
.C(n_5240),
.D(n_5246),
.Y(n_5302)
);

AOI22xp5_ASAP7_75t_L g5303 ( 
.A1(n_5265),
.A2(n_5244),
.B1(n_5226),
.B2(n_5233),
.Y(n_5303)
);

INVx1_ASAP7_75t_SL g5304 ( 
.A(n_5273),
.Y(n_5304)
);

AND3x4_ASAP7_75t_L g5305 ( 
.A(n_5258),
.B(n_5227),
.C(n_901),
.Y(n_5305)
);

NOR2xp67_ASAP7_75t_L g5306 ( 
.A(n_5264),
.B(n_5227),
.Y(n_5306)
);

NOR2x1_ASAP7_75t_L g5307 ( 
.A(n_5267),
.B(n_901),
.Y(n_5307)
);

INVxp67_ASAP7_75t_L g5308 ( 
.A(n_5281),
.Y(n_5308)
);

OAI221xp5_ASAP7_75t_L g5309 ( 
.A1(n_5292),
.A2(n_5266),
.B1(n_5282),
.B2(n_5278),
.C(n_5275),
.Y(n_5309)
);

OAI22xp33_ASAP7_75t_L g5310 ( 
.A1(n_5306),
.A2(n_5304),
.B1(n_5286),
.B2(n_5303),
.Y(n_5310)
);

AOI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_5301),
.A2(n_5269),
.B(n_5291),
.Y(n_5311)
);

OAI211xp5_ASAP7_75t_L g5312 ( 
.A1(n_5294),
.A2(n_5259),
.B(n_5287),
.C(n_5274),
.Y(n_5312)
);

OAI22xp5_ASAP7_75t_L g5313 ( 
.A1(n_5305),
.A2(n_5289),
.B1(n_5257),
.B2(n_5288),
.Y(n_5313)
);

NAND4xp25_ASAP7_75t_L g5314 ( 
.A(n_5300),
.B(n_5280),
.C(n_5272),
.D(n_5283),
.Y(n_5314)
);

OAI211xp5_ASAP7_75t_SL g5315 ( 
.A1(n_5308),
.A2(n_906),
.B(n_902),
.C(n_904),
.Y(n_5315)
);

NAND4xp25_ASAP7_75t_L g5316 ( 
.A(n_5295),
.B(n_906),
.C(n_902),
.D(n_904),
.Y(n_5316)
);

NAND4xp75_ASAP7_75t_L g5317 ( 
.A(n_5307),
.B(n_909),
.C(n_907),
.D(n_908),
.Y(n_5317)
);

OAI21xp5_ASAP7_75t_SL g5318 ( 
.A1(n_5297),
.A2(n_907),
.B(n_908),
.Y(n_5318)
);

AOI221xp5_ASAP7_75t_L g5319 ( 
.A1(n_5296),
.A2(n_912),
.B1(n_909),
.B2(n_910),
.C(n_913),
.Y(n_5319)
);

HB1xp67_ASAP7_75t_L g5320 ( 
.A(n_5317),
.Y(n_5320)
);

INVx3_ASAP7_75t_L g5321 ( 
.A(n_5315),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_L g5322 ( 
.A(n_5318),
.B(n_5316),
.Y(n_5322)
);

INVx3_ASAP7_75t_L g5323 ( 
.A(n_5310),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_5311),
.B(n_5293),
.Y(n_5324)
);

INVx2_ASAP7_75t_L g5325 ( 
.A(n_5309),
.Y(n_5325)
);

NAND3x1_ASAP7_75t_L g5326 ( 
.A(n_5319),
.B(n_5298),
.C(n_5299),
.Y(n_5326)
);

OR3x1_ASAP7_75t_L g5327 ( 
.A(n_5322),
.B(n_5314),
.C(n_5312),
.Y(n_5327)
);

INVx1_ASAP7_75t_SL g5328 ( 
.A(n_5320),
.Y(n_5328)
);

INVx5_ASAP7_75t_L g5329 ( 
.A(n_5323),
.Y(n_5329)
);

OR2x2_ASAP7_75t_L g5330 ( 
.A(n_5321),
.B(n_5313),
.Y(n_5330)
);

NOR2xp67_ASAP7_75t_L g5331 ( 
.A(n_5325),
.B(n_5324),
.Y(n_5331)
);

INVxp33_ASAP7_75t_SL g5332 ( 
.A(n_5328),
.Y(n_5332)
);

INVxp67_ASAP7_75t_L g5333 ( 
.A(n_5331),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5333),
.Y(n_5334)
);

INVxp67_ASAP7_75t_L g5335 ( 
.A(n_5334),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_5335),
.A2(n_5332),
.B(n_5330),
.Y(n_5336)
);

XNOR2xp5_ASAP7_75t_L g5337 ( 
.A(n_5336),
.B(n_5327),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_5337),
.B(n_5329),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_5338),
.A2(n_5302),
.B(n_5326),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5339),
.Y(n_5340)
);

AOI221xp5_ASAP7_75t_L g5341 ( 
.A1(n_5340),
.A2(n_913),
.B1(n_910),
.B2(n_912),
.C(n_914),
.Y(n_5341)
);

OR2x2_ASAP7_75t_L g5342 ( 
.A(n_5340),
.B(n_915),
.Y(n_5342)
);

AOI21xp5_ASAP7_75t_L g5343 ( 
.A1(n_5341),
.A2(n_916),
.B(n_917),
.Y(n_5343)
);

AOI211xp5_ASAP7_75t_L g5344 ( 
.A1(n_5343),
.A2(n_5342),
.B(n_919),
.C(n_917),
.Y(n_5344)
);


endmodule