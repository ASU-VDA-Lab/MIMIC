module fake_jpeg_25936_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_21),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_28),
.B(n_24),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_16),
.B(n_22),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.C(n_34),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_15),
.B1(n_27),
.B2(n_17),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_18),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_28),
.B(n_23),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_26),
.B1(n_13),
.B2(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_29),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_19),
.B(n_20),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.C(n_7),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_9),
.C(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);


endmodule