module fake_jpeg_506_n_80 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_21),
.B(n_19),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_26),
.B1(n_28),
.B2(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_40),
.B1(n_28),
.B2(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_29),
.B(n_27),
.C(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_38),
.B1(n_39),
.B2(n_37),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_54),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_56),
.B1(n_43),
.B2(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_23),
.B1(n_4),
.B2(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_63),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_17),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_3),
.C(n_4),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

OAI322xp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_59),
.C2(n_71),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_70),
.B1(n_63),
.B2(n_61),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_10),
.B(n_7),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_74),
.C(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_67),
.Y(n_76)
);

NOR2xp67_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_73),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_68),
.C(n_73),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_9),
.Y(n_80)
);


endmodule