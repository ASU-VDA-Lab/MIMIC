module fake_jpeg_18761_n_229 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_17),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_34),
.B(n_42),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_53),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_27),
.B1(n_11),
.B2(n_18),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_27),
.B1(n_11),
.B2(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_11),
.B1(n_28),
.B2(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_11),
.B1(n_24),
.B2(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_29),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_20),
.B1(n_21),
.B2(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_47),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_47),
.B(n_44),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_88),
.B(n_92),
.Y(n_109)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_71),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_47),
.C(n_49),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_68),
.C(n_67),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_48),
.B(n_38),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_48),
.B1(n_51),
.B2(n_29),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_96),
.B(n_72),
.C(n_41),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_17),
.B(n_13),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_65),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_43),
.B(n_29),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_110),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_82),
.C(n_86),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_70),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_13),
.B(n_17),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_65),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_38),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_117),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_85),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_81),
.B1(n_90),
.B2(n_84),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_97),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_124),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_94),
.B1(n_96),
.B2(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_82),
.B1(n_89),
.B2(n_86),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_141),
.B(n_13),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_94),
.B1(n_69),
.B2(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_131),
.B1(n_144),
.B2(n_50),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_142),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_139),
.C(n_116),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_113),
.B1(n_119),
.B2(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_90),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_90),
.C(n_84),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_117),
.B1(n_107),
.B2(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_16),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_154),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.C(n_160),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_116),
.C(n_45),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_23),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_135),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_133),
.C(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_127),
.B1(n_129),
.B2(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_162),
.B1(n_166),
.B2(n_172),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_131),
.B(n_128),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_172),
.B(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_125),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_131),
.B(n_138),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_52),
.C(n_79),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_149),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_191),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_156),
.C(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_79),
.C(n_41),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_160),
.C(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_188),
.Y(n_199)
);

NAND4xp25_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_23),
.C(n_52),
.D(n_45),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_189),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_158),
.C(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_177),
.B1(n_173),
.B2(n_57),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_177),
.B1(n_170),
.B2(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_200),
.B1(n_0),
.B2(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_168),
.B(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_31),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_186),
.B1(n_15),
.B2(n_16),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_23),
.B(n_7),
.Y(n_205)
);

AOI31xp67_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_209),
.A3(n_200),
.B(n_8),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_14),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_4),
.A3(n_9),
.B1(n_6),
.B2(n_5),
.C1(n_0),
.C2(n_3),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_31),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.C(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_5),
.Y(n_209)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_198),
.C(n_192),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_202),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_207),
.A2(n_30),
.B(n_5),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_4),
.B(n_6),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_220),
.B(n_1),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_4),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_0),
.C(n_1),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_211),
.B(n_9),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_222),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_224),
.C(n_219),
.Y(n_226)
);

BUFx12f_ASAP7_75t_SL g227 ( 
.A(n_226),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_225),
.B(n_2),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_2),
.Y(n_229)
);


endmodule