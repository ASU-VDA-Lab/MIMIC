module fake_netlist_6_1708_n_1131 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1131);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1131;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_209;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_1033;
wire n_208;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_168;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_953;
wire n_1017;
wire n_1004;
wire n_448;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_689;
wire n_231;
wire n_354;
wire n_409;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_195;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_834;
wire n_207;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_165;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_170;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_169;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_93),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_76),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_62),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_55),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_28),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_84),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_58),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_49),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_43),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_79),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_48),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_4),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_68),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_122),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_34),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_57),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_50),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_123),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_17),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_125),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_60),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_88),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_159),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_67),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_172),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_175),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_194),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_232),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx12_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_228),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_225),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_226),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_233),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_220),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_234),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_232),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_218),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_218),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_244),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_218),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_232),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_218),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_218),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_272),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_204),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_294),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_272),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_292),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_269),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_269),
.Y(n_322)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_250),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_277),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_258),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_266),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_338),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_249),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_315),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_253),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_338),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_310),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_296),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_323),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_306),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_315),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_322),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_253),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_321),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_326),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_321),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_337),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_339),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_342),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_339),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_254),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_383),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_346),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_267),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_374),
.B(n_179),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_361),
.B(n_179),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

CKINVDCx11_ASAP7_75t_R g404 ( 
.A(n_343),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_331),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_369),
.A2(n_312),
.B(n_300),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_349),
.B(n_192),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_328),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_344),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_329),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_373),
.B(n_299),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_387),
.A2(n_301),
.B(n_320),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_353),
.B(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g426 ( 
.A(n_355),
.B(n_326),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_335),
.Y(n_427)
);

BUFx8_ASAP7_75t_SL g428 ( 
.A(n_343),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_359),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_387),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_371),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_350),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_L g438 ( 
.A1(n_366),
.A2(n_341),
.B1(n_340),
.B2(n_163),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_366),
.Y(n_439)
);

NOR2x1_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_340),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_344),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_343),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_374),
.B(n_192),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_345),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_385),
.B(n_341),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_345),
.B(n_309),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_358),
.A2(n_327),
.B(n_324),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_345),
.B(n_268),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_345),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_345),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_345),
.B(n_273),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_362),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_345),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_345),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_374),
.B(n_200),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_345),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_345),
.B(n_286),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_343),
.Y(n_470)
);

AOI22x1_ASAP7_75t_SL g471 ( 
.A1(n_343),
.A2(n_210),
.B1(n_191),
.B2(n_196),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_396),
.B(n_254),
.Y(n_473)
);

NAND2x1_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_326),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_390),
.B(n_287),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_418),
.B(n_290),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_415),
.A2(n_210),
.B1(n_200),
.B2(n_167),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_295),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_396),
.B(n_274),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_415),
.A2(n_274),
.B1(n_293),
.B2(n_291),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_401),
.B(n_447),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_403),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g496 ( 
.A(n_418),
.B(n_291),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_397),
.B(n_293),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_182),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_447),
.B(n_326),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_401),
.B(n_170),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_397),
.B(n_326),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_390),
.B(n_187),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_458),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_416),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_197),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_457),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_464),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_486),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_486),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_486),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_416),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_424),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_486),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_488),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_492),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_488),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_477),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_484),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_481),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_482),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_495),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_517),
.A2(n_410),
.B(n_423),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_514),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_514),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_476),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_475),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_483),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_473),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_479),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_R g546 ( 
.A(n_497),
.B(n_441),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_491),
.B(n_422),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_518),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_R g550 ( 
.A(n_485),
.B(n_441),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_507),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_485),
.B(n_419),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_507),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_507),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_501),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_525),
.B(n_487),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_487),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_480),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_548),
.A2(n_480),
.B1(n_493),
.B2(n_438),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_528),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_489),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_530),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_535),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_536),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_541),
.B(n_429),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_392),
.C(n_500),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_537),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_500),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_552),
.B(n_493),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_539),
.B(n_489),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_545),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_540),
.B(n_439),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_521),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_538),
.Y(n_583)
);

AND3x2_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_392),
.C(n_511),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_511),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_544),
.B(n_424),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_SL g589 ( 
.A1(n_547),
.A2(n_493),
.B(n_499),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_538),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_532),
.B(n_459),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_547),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_538),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_527),
.A2(n_438),
.B1(n_407),
.B2(n_425),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_524),
.A2(n_436),
.B1(n_432),
.B2(n_434),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_528),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_528),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_526),
.B(n_435),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_525),
.A2(n_407),
.B1(n_430),
.B2(n_501),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_526),
.B(n_459),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_R g609 ( 
.A(n_550),
.B(n_429),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_526),
.B(n_469),
.C(n_462),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_528),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_548),
.A2(n_471),
.B1(n_517),
.B2(n_512),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_528),
.B(n_404),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_526),
.A2(n_503),
.B1(n_506),
.B2(n_502),
.Y(n_614)
);

INVx6_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_520),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_526),
.B(n_433),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_554),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_526),
.B(n_462),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_533),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_526),
.A2(n_503),
.B1(n_506),
.B2(n_502),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_531),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_469),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_526),
.B(n_505),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_521),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_531),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_585),
.B(n_426),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_443),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_618),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_606),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_596),
.B(n_435),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_558),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_626),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_564),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_560),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_588),
.B(n_428),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_577),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_597),
.B(n_508),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_605),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_563),
.A2(n_516),
.B1(n_509),
.B2(n_513),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_610),
.B(n_419),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_580),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_613),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_562),
.B(n_412),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_575),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_572),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_595),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_618),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_573),
.B(n_428),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_616),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_563),
.B(n_419),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_570),
.B(n_419),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_555),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_559),
.B(n_516),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_567),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_627),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_555),
.B(n_508),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_628),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_591),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_604),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_605),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_617),
.B(n_420),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_611),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_581),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_579),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_581),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_440),
.C(n_398),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_582),
.B(n_509),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_557),
.B(n_513),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_557),
.B(n_490),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_586),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_623),
.B(n_417),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_556),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_576),
.B(n_594),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_607),
.B(n_614),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_576),
.B(n_494),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_599),
.B(n_431),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_574),
.B(n_474),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_613),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_607),
.B(n_515),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_614),
.B(n_478),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_581),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_594),
.B(n_620),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_574),
.B(n_498),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_581),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_608),
.B(n_470),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_568),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_625),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_619),
.B(n_624),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_625),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_625),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_617),
.B(n_453),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_652),
.B(n_624),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_636),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_682),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_638),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_631),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_671),
.B(n_619),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_690),
.B(n_687),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_660),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_689),
.B(n_584),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_631),
.Y(n_716)
);

OAI221xp5_ASAP7_75t_L g717 ( 
.A1(n_689),
.A2(n_621),
.B1(n_603),
.B2(n_569),
.C(n_589),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_664),
.B(n_598),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_667),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_656),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_683),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_670),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_701),
.B(n_584),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_685),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_640),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_671),
.B(n_601),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_655),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_634),
.B(n_621),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_657),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_695),
.B(n_620),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_695),
.B(n_587),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_641),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_664),
.B(n_598),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_675),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_663),
.B(n_601),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_662),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_634),
.B(n_592),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_675),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_666),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_677),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_699),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_656),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_635),
.B(n_612),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_645),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_661),
.A2(n_612),
.B1(n_600),
.B2(n_467),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_648),
.B(n_578),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_692),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_687),
.A2(n_590),
.B1(n_593),
.B2(n_583),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_656),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_662),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_637),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_653),
.B(n_417),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_680),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_650),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_668),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_669),
.B(n_625),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_680),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_669),
.B(n_602),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_653),
.B(n_583),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_692),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_668),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_677),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_632),
.B(n_602),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_674),
.A2(n_612),
.B1(n_609),
.B2(n_453),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_691),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_767),
.A2(n_698),
.B1(n_684),
.B2(n_696),
.C(n_630),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_708),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_742),
.B(n_765),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_715),
.A2(n_679),
.B1(n_609),
.B2(n_642),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_711),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_768),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_765),
.B(n_665),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_711),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_706),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_715),
.A2(n_679),
.B1(n_704),
.B2(n_647),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_723),
.A2(n_647),
.B1(n_629),
.B2(n_639),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_723),
.B(n_632),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_718),
.B(n_672),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_710),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_747),
.B(n_633),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_717),
.A2(n_693),
.B(n_498),
.C(n_450),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_726),
.B(n_633),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_721),
.B(n_646),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_724),
.B(n_690),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_717),
.A2(n_467),
.B1(n_690),
.B2(n_404),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_SL g789 ( 
.A(n_707),
.B(n_646),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_737),
.B(n_673),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_766),
.B(n_673),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_714),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_766),
.B(n_681),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_761),
.B(n_643),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_749),
.B(n_686),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_719),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_722),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_737),
.B(n_393),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_749),
.B(n_686),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_735),
.B(n_651),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_729),
.B(n_411),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_761),
.B(n_643),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_712),
.B(n_686),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_707),
.B(n_644),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_713),
.A2(n_745),
.B1(n_705),
.B2(n_747),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_755),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_713),
.A2(n_467),
.B1(n_186),
.B2(n_209),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_707),
.A2(n_644),
.B(n_593),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_707),
.B(n_649),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_757),
.B(n_649),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_713),
.B(n_697),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_711),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_727),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_730),
.B(n_668),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_763),
.B(n_721),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_728),
.B(n_590),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_730),
.B(n_678),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_709),
.B(n_697),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_736),
.B(n_678),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_728),
.B(n_651),
.Y(n_821)
);

AND2x6_ASAP7_75t_SL g822 ( 
.A(n_748),
.B(n_395),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_739),
.B(n_676),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_740),
.A2(n_615),
.B1(n_450),
.B2(n_463),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_716),
.B(n_678),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_762),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_716),
.B(n_744),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_756),
.B(n_676),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_729),
.B(n_466),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_720),
.B(n_395),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_754),
.B(n_700),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_760),
.B(n_703),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_744),
.B(n_412),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_732),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_771),
.B(n_746),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_786),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_789),
.B(n_751),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_806),
.B(n_751),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_811),
.B(n_731),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_817),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_821),
.B(n_750),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_775),
.B(n_725),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_786),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_780),
.B(n_751),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_782),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_792),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_797),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_774),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_790),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_781),
.Y(n_851)
);

AND2x2_ASAP7_75t_SL g852 ( 
.A(n_783),
.B(n_759),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_796),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_784),
.A2(n_772),
.B(n_788),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_811),
.B(n_731),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_800),
.B(n_733),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_795),
.B(n_734),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_826),
.B(n_813),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_834),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_770),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_819),
.B(n_741),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_819),
.B(n_743),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_815),
.Y(n_863)
);

BUFx4f_ASAP7_75t_L g864 ( 
.A(n_817),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_809),
.B(n_738),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_785),
.B(n_738),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_817),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_810),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_831),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_808),
.B(n_644),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_828),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_803),
.B(n_769),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_828),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_827),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_823),
.B(n_758),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_787),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_799),
.B(n_764),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_822),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_804),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_816),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_832),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_863),
.B(n_881),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_854),
.A2(n_791),
.B(n_793),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_849),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_852),
.A2(n_805),
.B1(n_778),
.B2(n_779),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_852),
.A2(n_802),
.B(n_794),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_869),
.B(n_842),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_874),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_801),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_869),
.B(n_876),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_857),
.A2(n_798),
.B(n_814),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_857),
.A2(n_818),
.B(n_807),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_872),
.A2(n_829),
.B(n_820),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_872),
.A2(n_824),
.B(n_830),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_850),
.A2(n_825),
.B(n_833),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_874),
.B(n_752),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_879),
.B(n_773),
.Y(n_898)
);

AO21x1_ASAP7_75t_L g899 ( 
.A1(n_879),
.A2(n_202),
.B(n_201),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_850),
.A2(n_812),
.B(n_776),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_837),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_870),
.A2(n_463),
.B(n_703),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_836),
.B(n_827),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_846),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_870),
.A2(n_688),
.B(n_682),
.Y(n_905)
);

OAI321xp33_ASAP7_75t_L g906 ( 
.A1(n_838),
.A2(n_180),
.A3(n_186),
.B1(n_209),
.B2(n_214),
.C(n_764),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_868),
.A2(n_186),
.B(n_209),
.C(n_180),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_849),
.B(n_764),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_871),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_871),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_840),
.A2(n_622),
.B(n_753),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_843),
.A2(n_186),
.B(n_180),
.Y(n_913)
);

NAND2x1_ASAP7_75t_L g914 ( 
.A(n_836),
.B(n_682),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_858),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_845),
.A2(n_180),
.B(n_209),
.C(n_214),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_839),
.A2(n_214),
.B(n_198),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_841),
.B(n_694),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_844),
.B(n_694),
.Y(n_919)
);

AO21x1_ASAP7_75t_L g920 ( 
.A1(n_841),
.A2(n_0),
.B(n_1),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_880),
.B(n_702),
.Y(n_921)
);

AOI33xp33_ASAP7_75t_L g922 ( 
.A1(n_859),
.A2(n_421),
.A3(n_408),
.B1(n_409),
.B2(n_3),
.B3(n_4),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_851),
.B(n_0),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_855),
.A2(n_864),
.B(n_878),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_899),
.A2(n_864),
.B(n_855),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_903),
.B(n_844),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_922),
.A2(n_855),
.B(n_865),
.C(n_880),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_916),
.A2(n_867),
.B(n_860),
.C(n_865),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_886),
.A2(n_880),
.B(n_847),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_884),
.A2(n_880),
.B(n_847),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_895),
.A2(n_860),
.B(n_861),
.Y(n_931)
);

CKINVDCx8_ASAP7_75t_R g932 ( 
.A(n_897),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_896),
.B(n_856),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_883),
.B(n_875),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_888),
.B(n_848),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_907),
.A2(n_862),
.B(n_866),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_910),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_913),
.A2(n_835),
.B(n_848),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_913),
.A2(n_882),
.B1(n_877),
.B2(n_873),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_892),
.B(n_871),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_890),
.B(n_873),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_894),
.A2(n_841),
.B(n_867),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_932),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_929),
.A2(n_920),
.B(n_902),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_942),
.B(n_889),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_SL g946 ( 
.A1(n_942),
.A2(n_885),
.B1(n_923),
.B2(n_898),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_930),
.A2(n_900),
.B(n_915),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_927),
.B(n_889),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_933),
.B(n_908),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_935),
.B(n_891),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_925),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_931),
.B(n_887),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_928),
.A2(n_917),
.B(n_893),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_926),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_940),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_941),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_934),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_939),
.Y(n_959)
);

CKINVDCx14_ASAP7_75t_R g960 ( 
.A(n_936),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_938),
.B(n_901),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_927),
.B(n_904),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_929),
.A2(n_906),
.B(n_924),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_932),
.B(n_1),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_935),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_926),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_965),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_945),
.B(n_919),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_945),
.B(n_910),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_967),
.B(n_909),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_961),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_952),
.B(n_944),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_960),
.A2(n_905),
.B(n_914),
.C(n_912),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_958),
.B(n_911),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_973),
.A2(n_953),
.B(n_954),
.C(n_963),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_972),
.B(n_962),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_977),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_976),
.A2(n_946),
.B(n_949),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_979),
.A2(n_948),
.B(n_947),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_978),
.B(n_968),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_980),
.A2(n_948),
.B(n_947),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_981),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_983),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_982),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_985),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_984),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_987),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_986),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_986),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_988),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_989),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_991),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_992),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_995),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_995),
.B(n_984),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_997),
.B(n_993),
.Y(n_998)
);

INVx5_ASAP7_75t_SL g999 ( 
.A(n_996),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_998),
.B(n_994),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_999),
.Y(n_1001)
);

NAND2x1_ASAP7_75t_L g1002 ( 
.A(n_1000),
.B(n_943),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_1001),
.B(n_970),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1002),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_1003),
.B(n_969),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_1005),
.B(n_982),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_957),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_1005),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1006),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_1007),
.B(n_957),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1008),
.B(n_957),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1011),
.B(n_1010),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_1009),
.B(n_943),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_1013),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1012),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_966),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1015),
.B(n_943),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1017),
.B(n_956),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1019),
.B(n_956),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_1021),
.B(n_956),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1020),
.Y(n_1023)
);

OAI22xp33_ASAP7_75t_SL g1024 ( 
.A1(n_1023),
.A2(n_421),
.B1(n_959),
.B2(n_199),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_1022),
.A2(n_975),
.B1(n_955),
.B2(n_950),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_2),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1024),
.B(n_2),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1027),
.A2(n_203),
.B(n_195),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1030),
.B(n_1029),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1031),
.B(n_3),
.Y(n_1033)
);

XNOR2x2_ASAP7_75t_SL g1034 ( 
.A(n_1032),
.B(n_206),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1033),
.B(n_970),
.Y(n_1035)
);

AOI32xp33_ASAP7_75t_L g1036 ( 
.A1(n_1035),
.A2(n_212),
.A3(n_208),
.B1(n_211),
.B2(n_213),
.Y(n_1036)
);

AOI222xp33_ASAP7_75t_L g1037 ( 
.A1(n_1034),
.A2(n_214),
.B1(n_207),
.B2(n_975),
.C1(n_974),
.C2(n_467),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1036),
.Y(n_1038)
);

AOI211x1_ASAP7_75t_L g1039 ( 
.A1(n_1037),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1038),
.Y(n_1040)
);

AOI31xp33_ASAP7_75t_L g1041 ( 
.A1(n_1039),
.A2(n_964),
.A3(n_7),
.B(n_8),
.Y(n_1041)
);

NAND5xp2_ASAP7_75t_L g1042 ( 
.A(n_1040),
.B(n_6),
.C(n_9),
.D(n_10),
.E(n_11),
.Y(n_1042)
);

AOI211xp5_ASAP7_75t_SL g1043 ( 
.A1(n_1041),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_1040),
.B(n_12),
.C(n_13),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1042),
.B(n_12),
.Y(n_1045)
);

OAI221xp5_ASAP7_75t_SL g1046 ( 
.A1(n_1043),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_1046)
);

OAI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1044),
.A2(n_389),
.B1(n_445),
.B2(n_448),
.Y(n_1047)
);

NAND4xp25_ASAP7_75t_SL g1048 ( 
.A(n_1045),
.B(n_14),
.C(n_16),
.D(n_17),
.Y(n_1048)
);

NAND5xp2_ASAP7_75t_L g1049 ( 
.A(n_1046),
.B(n_18),
.C(n_19),
.D(n_20),
.E(n_21),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_1049),
.B(n_1047),
.C(n_18),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1048),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_445),
.B1(n_448),
.B2(n_449),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_19),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_1053),
.B(n_21),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_SL g1055 ( 
.A(n_1052),
.B(n_445),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1055),
.B(n_448),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_449),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_1056),
.B(n_22),
.Y(n_1058)
);

NOR4xp75_ASAP7_75t_L g1059 ( 
.A(n_1057),
.B(n_22),
.C(n_23),
.D(n_24),
.Y(n_1059)
);

XOR2x1_ASAP7_75t_L g1060 ( 
.A(n_1059),
.B(n_23),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1058),
.B(n_24),
.C(n_25),
.Y(n_1061)
);

AOI211xp5_ASAP7_75t_L g1062 ( 
.A1(n_1058),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1062)
);

XNOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1060),
.B(n_26),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_1061),
.Y(n_1064)
);

NAND4xp75_ASAP7_75t_L g1065 ( 
.A(n_1062),
.B(n_27),
.C(n_28),
.D(n_29),
.Y(n_1065)
);

AO22x2_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1066)
);

AO22x2_ASAP7_75t_L g1067 ( 
.A1(n_1063),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1067),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1066),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1069),
.B(n_1065),
.Y(n_1070)
);

OA22x2_ASAP7_75t_L g1071 ( 
.A1(n_1068),
.A2(n_971),
.B1(n_38),
.B2(n_39),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1070),
.A2(n_472),
.B1(n_449),
.B2(n_406),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1071),
.Y(n_1073)
);

OAI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1073),
.A2(n_472),
.B1(n_40),
.B2(n_41),
.C(n_42),
.Y(n_1074)
);

NAND5xp2_ASAP7_75t_L g1075 ( 
.A(n_1072),
.B(n_37),
.C(n_44),
.D(n_45),
.E(n_46),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1074),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1076),
.A2(n_472),
.B1(n_406),
.B2(n_897),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_406),
.B1(n_897),
.B2(n_468),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_1076),
.A2(n_47),
.B(n_51),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1079),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1078),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

AO22x1_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1085)
);

OAI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1082),
.A2(n_951),
.B1(n_59),
.B2(n_61),
.C1(n_65),
.C2(n_69),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1084),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_1085),
.B(n_56),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1086),
.Y(n_1089)
);

AOI222xp33_ASAP7_75t_L g1090 ( 
.A1(n_1087),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C1(n_73),
.C2(n_74),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1089),
.Y(n_1091)
);

OAI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1088),
.A2(n_398),
.B1(n_397),
.B2(n_918),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1091),
.A2(n_897),
.B(n_921),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1092),
.A2(n_75),
.B(n_77),
.Y(n_1094)
);

AO221x2_ASAP7_75t_L g1095 ( 
.A1(n_1090),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.C(n_82),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1091),
.B(n_83),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1091),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1091),
.A2(n_398),
.B1(n_504),
.B2(n_89),
.Y(n_1098)
);

AOI211xp5_ASAP7_75t_L g1099 ( 
.A1(n_1091),
.A2(n_85),
.B(n_87),
.C(n_90),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1091),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1091),
.A2(n_92),
.B(n_95),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1091),
.B(n_96),
.Y(n_1102)
);

OAI211xp5_ASAP7_75t_L g1103 ( 
.A1(n_1091),
.A2(n_97),
.B(n_100),
.C(n_101),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1091),
.A2(n_103),
.B(n_104),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1091),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1100),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1105),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1097),
.B(n_105),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1094),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1095),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1095),
.Y(n_1111)
);

OR3x1_ASAP7_75t_L g1112 ( 
.A(n_1102),
.B(n_106),
.C(n_107),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1096),
.A2(n_504),
.B1(n_110),
.B2(n_111),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1104),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1106),
.A2(n_1098),
.B1(n_1103),
.B2(n_1101),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1093),
.B2(n_615),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1109),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_R g1118 ( 
.A1(n_1114),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_1110),
.A2(n_118),
.B(n_119),
.Y(n_1119)
);

AOI222xp33_ASAP7_75t_L g1120 ( 
.A1(n_1111),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.C1(n_126),
.C2(n_127),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1115),
.A2(n_1112),
.B(n_1113),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1116),
.B(n_1108),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1119),
.B(n_128),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_1117),
.B1(n_1118),
.B2(n_1120),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_1121),
.B1(n_1123),
.B2(n_136),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1125),
.B(n_131),
.Y(n_1126)
);

OAI221xp5_ASAP7_75t_R g1127 ( 
.A1(n_1126),
.A2(n_133),
.B1(n_138),
.B2(n_139),
.C(n_140),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1127),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.C(n_145),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1128),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_1129)
);

AOI211xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1130)
);

AOI211xp5_ASAP7_75t_L g1131 ( 
.A1(n_1130),
.A2(n_153),
.B(n_154),
.C(n_156),
.Y(n_1131)
);


endmodule