module real_jpeg_15526_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_216;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_1),
.Y(n_138)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_4),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_40),
.B1(n_61),
.B2(n_65),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_7),
.B(n_85),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_136),
.C(n_139),
.Y(n_135)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_168),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI21x1_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_126),
.B(n_167),
.Y(n_11)
);

NOR2xp67_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_121),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_13),
.B(n_121),
.Y(n_167)
);

XOR2x2_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_82),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_58),
.B2(n_59),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_15),
.B(n_82),
.C(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_17),
.B(n_124),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.A3(n_26),
.B1(n_32),
.B2(n_36),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_35),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_36),
.A2(n_40),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_40),
.B(n_69),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_40),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_40),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_40),
.A2(n_204),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_41),
.A2(n_42),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_41),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_41),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_41),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_41),
.A2(n_124),
.B1(n_177),
.B2(n_207),
.Y(n_176)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_83),
.B(n_122),
.C(n_125),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_59),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_59),
.B1(n_134),
.B2(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_58),
.B(n_124),
.C(n_132),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_58),
.A2(n_59),
.B1(n_83),
.B2(n_120),
.Y(n_165)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_84),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_87),
.B1(n_90),
.B2(n_92),
.Y(n_86)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_108),
.B1(n_119),
.B2(n_120),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_83),
.B(n_110),
.C(n_124),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B(n_105),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_112),
.B(n_217),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_123),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_130),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_161),
.B(n_166),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_142),
.B(n_160),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_133),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_157),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_222),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_173),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_208),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_193),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_198),
.B(n_203),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);


endmodule