module real_jpeg_3768_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_66),
.B1(n_74),
.B2(n_101),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_1),
.A2(n_66),
.B1(n_129),
.B2(n_277),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_1),
.A2(n_66),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_73),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_3),
.A2(n_73),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_73),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_3),
.B(n_90),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_258),
.B(n_260),
.C(n_264),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_3),
.B(n_289),
.C(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_3),
.B(n_69),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_3),
.B(n_114),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_6),
.Y(n_316)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_6),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_10),
.Y(n_169)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_10),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_10),
.Y(n_182)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_12),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_58),
.B1(n_140),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_12),
.A2(n_58),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_58),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_13),
.A2(n_134),
.B1(n_135),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_134),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_230),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_228),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_195),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_22),
.B(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_22),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_22),
.B(n_232),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_131),
.CI(n_158),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_70),
.C(n_102),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_24),
.A2(n_102),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_24),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_61),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_53),
.Y(n_26)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_43),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_35),
.Y(n_266)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_36),
.Y(n_166)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_42),
.Y(n_192)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_43),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_47),
.Y(n_157)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_47),
.Y(n_218)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_52),
.Y(n_259)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_54),
.B(n_69),
.Y(n_241)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_61),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_62),
.B(n_194),
.Y(n_193)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_69),
.A2(n_188),
.B(n_194),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_70),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_99),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_73),
.A2(n_261),
.B(n_263),
.Y(n_260)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_78),
.B(n_100),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_78),
.B(n_178),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_90),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_178),
.Y(n_177)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_99),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_102),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_123),
.B(n_124),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_104),
.B(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_104),
.B(n_276),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_105)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_115),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_114),
.B(n_276),
.Y(n_293)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_118),
.Y(n_302)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_122),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_122),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_123),
.A2(n_212),
.B(n_219),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_123),
.B(n_124),
.Y(n_274)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_128),
.Y(n_287)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_150),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_132),
.B(n_150),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_142),
.B(n_147),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_143),
.B(n_204),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_143),
.A2(n_204),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_143),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_147),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_147),
.B(n_297),
.Y(n_327)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_151),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_152),
.B(n_275),
.Y(n_304)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_176),
.C(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_164),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.A3(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_188),
.B(n_194),
.Y(n_339)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_220),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_211),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_200),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_207),
.Y(n_301)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_210),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_219),
.B(n_293),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_246),
.B(n_351),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_239),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_245),
.B(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_280),
.B(n_350),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_249),
.B(n_252),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_271),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_256),
.A2(n_271),
.B1(n_272),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_256),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_267),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_257),
.A2(n_267),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_344),
.B(n_349),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_332),
.B(n_343),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_308),
.B(n_331),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_286),
.B1(n_292),
.B2(n_311),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_306),
.C(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_317),
.B(n_330),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_312),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_326),
.B(n_329),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_335),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.C(n_340),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_348),
.Y(n_349)
);


endmodule