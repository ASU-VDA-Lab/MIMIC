module fake_jpeg_14096_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_62),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_66),
.Y(n_222)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_68),
.B(n_69),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_20),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_74),
.B(n_76),
.Y(n_162)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_86),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_20),
.B(n_16),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_90),
.B(n_94),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_93),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_15),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_96),
.B(n_97),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_99),
.B(n_103),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_100),
.A2(n_40),
.B1(n_46),
.B2(n_41),
.Y(n_216)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_0),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_47),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_111),
.B(n_112),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_48),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_0),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_126),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_48),
.B(n_0),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_40),
.Y(n_137)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_137),
.B(n_175),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

BUFx4f_ASAP7_75t_SL g259 ( 
.A(n_138),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_140),
.B(n_184),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_145),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_64),
.A2(n_83),
.B(n_106),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_152),
.B(n_30),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_59),
.B(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_217),
.Y(n_223)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_107),
.A2(n_51),
.B1(n_56),
.B2(n_28),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_179),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_181),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_65),
.B(n_27),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_75),
.B(n_82),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_12),
.Y(n_275)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_66),
.A2(n_53),
.B1(n_55),
.B2(n_30),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_218),
.B1(n_105),
.B2(n_95),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_67),
.B(n_27),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_203),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_81),
.B(n_55),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_195),
.B(n_139),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_60),
.Y(n_200)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_26),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_129),
.B(n_26),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_33),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_33),
.B1(n_41),
.B2(n_36),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_118),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_120),
.A2(n_53),
.B1(n_21),
.B2(n_23),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_227),
.A2(n_254),
.B1(n_210),
.B2(n_168),
.Y(n_317)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_228),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_132),
.A2(n_119),
.B1(n_114),
.B2(n_104),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_230),
.A2(n_235),
.B1(n_248),
.B2(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_146),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_231),
.B(n_241),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_232),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_195),
.B1(n_80),
.B2(n_88),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_233),
.A2(n_273),
.B1(n_173),
.B2(n_142),
.Y(n_329)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_183),
.A2(n_73),
.B1(n_72),
.B2(n_89),
.Y(n_235)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_21),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_242),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_105),
.B1(n_95),
.B2(n_23),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_243),
.A2(n_249),
.B(n_268),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_161),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_77),
.B1(n_29),
.B2(n_34),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_250),
.B(n_263),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_251),
.A2(n_258),
.B1(n_264),
.B2(n_198),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_253),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_157),
.A2(n_28),
.B1(n_34),
.B2(n_29),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_257),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_36),
.B1(n_2),
.B2(n_4),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_189),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_202),
.B(n_6),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_222),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_162),
.B(n_9),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_265),
.B(n_269),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_161),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_267),
.B(n_278),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_268),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_162),
.B(n_9),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_180),
.Y(n_270)
);

NAND2xp67_ASAP7_75t_SL g357 ( 
.A(n_270),
.B(n_289),
.Y(n_357)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_156),
.B(n_10),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_274),
.B(n_277),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_294),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_156),
.B(n_13),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_176),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_170),
.A2(n_13),
.B1(n_176),
.B2(n_218),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_261),
.B1(n_266),
.B2(n_239),
.Y(n_356)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_196),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_286),
.Y(n_305)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_154),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_163),
.B(n_190),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_138),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_288),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_208),
.B(n_169),
.Y(n_288)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_136),
.Y(n_290)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_133),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_199),
.B(n_155),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_293),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_153),
.B(n_185),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_164),
.B(n_148),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_196),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_295),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_135),
.Y(n_296)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_144),
.B(n_130),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_134),
.B(n_136),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_182),
.Y(n_300)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_177),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_301),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_235),
.A2(n_198),
.B1(n_173),
.B2(n_142),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_303),
.A2(n_356),
.B1(n_258),
.B2(n_291),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_317),
.B(n_245),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_229),
.B(n_171),
.C(n_210),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_321),
.B(n_322),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_249),
.B(n_135),
.C(n_174),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_237),
.B(n_166),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_341),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_225),
.B(n_215),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_327),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_346),
.B1(n_280),
.B2(n_255),
.Y(n_364)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_270),
.A2(n_194),
.B1(n_205),
.B2(n_201),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_333),
.A2(n_335),
.B1(n_343),
.B2(n_245),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_275),
.B(n_221),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_337),
.B(n_228),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_240),
.A2(n_200),
.B1(n_145),
.B2(n_181),
.Y(n_335)
);

AOI22x1_ASAP7_75t_L g337 ( 
.A1(n_275),
.A2(n_174),
.B1(n_149),
.B2(n_159),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_223),
.B(n_149),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_251),
.A2(n_204),
.B1(n_159),
.B2(n_165),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_273),
.A2(n_165),
.B1(n_193),
.B2(n_141),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_345),
.A2(n_266),
.B1(n_239),
.B2(n_272),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_243),
.A2(n_193),
.B1(n_219),
.B2(n_241),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_264),
.Y(n_362)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_247),
.Y(n_349)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

AND2x2_ASAP7_75t_SL g351 ( 
.A(n_294),
.B(n_260),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_351),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_262),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_352),
.B(n_246),
.Y(n_392)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_256),
.B(n_271),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_360),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_362),
.A2(n_367),
.B(n_370),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_364),
.A2(n_328),
.B1(n_356),
.B2(n_317),
.Y(n_410)
);

INVx11_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_236),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_366),
.B(n_373),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_259),
.Y(n_371)
);

AOI31xp33_ASAP7_75t_SL g442 ( 
.A1(n_371),
.A2(n_405),
.A3(n_398),
.B(n_367),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_285),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

CKINVDCx10_ASAP7_75t_R g376 ( 
.A(n_323),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_376),
.Y(n_438)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_348),
.A2(n_244),
.B(n_224),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_384),
.B(n_391),
.Y(n_413)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_315),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_386),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_283),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_385),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_224),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_320),
.B(n_234),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_399),
.Y(n_426)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_392),
.B(n_307),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_311),
.B(n_244),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_401),
.Y(n_441)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_395),
.Y(n_411)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_396),
.Y(n_421)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_397),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_302),
.B(n_246),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_300),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_259),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_312),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_290),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_404),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_259),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_238),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_328),
.A2(n_232),
.B1(n_253),
.B2(n_257),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_407),
.Y(n_429)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_322),
.B(n_296),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_360),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_410),
.A2(n_387),
.B1(n_365),
.B2(n_382),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_351),
.B(n_357),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_437),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_413),
.A2(n_437),
.B(n_375),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_415),
.B(n_418),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_368),
.A2(n_351),
.B1(n_321),
.B2(n_337),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_416),
.A2(n_430),
.B1(n_433),
.B2(n_434),
.Y(n_456)
);

XOR2x1_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_372),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_352),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_427),
.C(n_440),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_366),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_424),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_388),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_376),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_238),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_327),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_370),
.A2(n_337),
.B1(n_355),
.B2(n_327),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_363),
.A2(n_346),
.B1(n_307),
.B2(n_342),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_363),
.A2(n_307),
.B1(n_334),
.B2(n_316),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_424),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_380),
.A2(n_326),
.B(n_361),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_312),
.Y(n_440)
);

INVx6_ASAP7_75t_SL g449 ( 
.A(n_442),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_385),
.C(n_373),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_318),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_383),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_451),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_445),
.Y(n_451)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_453),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_435),
.A2(n_364),
.B1(n_403),
.B2(n_386),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_457),
.B1(n_472),
.B2(n_482),
.Y(n_487)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_455),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_435),
.A2(n_404),
.B1(n_406),
.B2(n_405),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_410),
.A2(n_369),
.B1(n_387),
.B2(n_407),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_477),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_461),
.B(n_444),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_462),
.A2(n_478),
.B(n_413),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_393),
.Y(n_463)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_371),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_SL g498 ( 
.A(n_464),
.B(n_430),
.C(n_417),
.Y(n_498)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_414),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_467),
.B(n_473),
.Y(n_494)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_469),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_414),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_433),
.C(n_434),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_471),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_429),
.A2(n_374),
.B1(n_378),
.B2(n_390),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_426),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_446),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_474),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_393),
.Y(n_475)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_475),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_476),
.A2(n_417),
.B(n_412),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_429),
.A2(n_441),
.B1(n_409),
.B2(n_420),
.Y(n_477)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_428),
.B(n_390),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_479),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_428),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_480),
.Y(n_511)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_411),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_436),
.A2(n_378),
.B1(n_374),
.B2(n_379),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_411),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_483),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_418),
.C(n_419),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_484),
.B(n_497),
.C(n_508),
.Y(n_534)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_491),
.A2(n_498),
.B(n_501),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_440),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_503),
.Y(n_526)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_496),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_415),
.C(n_427),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_499),
.B(n_497),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_500),
.B(n_510),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_478),
.A2(n_416),
.B(n_425),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_379),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_438),
.C(n_439),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_456),
.B(n_453),
.C(n_478),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_513),
.C(n_481),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_449),
.A2(n_448),
.B(n_476),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_456),
.B(n_479),
.C(n_463),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_432),
.B(n_421),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_421),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_496),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_518),
.B(n_529),
.Y(n_552)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_515),
.Y(n_520)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_520),
.Y(n_554)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_515),
.Y(n_521)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

BUFx5_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_479),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_527),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_524),
.B(n_486),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_489),
.A2(n_511),
.B1(n_490),
.B2(n_487),
.Y(n_525)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_525),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_484),
.B(n_475),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_490),
.A2(n_460),
.B1(n_464),
.B2(n_457),
.Y(n_528)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_528),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_494),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_517),
.A2(n_454),
.B1(n_472),
.B2(n_482),
.Y(n_530)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_532),
.A2(n_547),
.B(n_502),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_397),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_533),
.B(n_543),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_517),
.A2(n_493),
.B1(n_509),
.B2(n_513),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_538),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_491),
.Y(n_559)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_493),
.B(n_466),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_537),
.B(n_540),
.Y(n_561)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_512),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_495),
.A2(n_465),
.B1(n_458),
.B2(n_455),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_539),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_487),
.A2(n_469),
.B1(n_468),
.B2(n_439),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_541),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_512),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_544),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_502),
.A2(n_432),
.B1(n_377),
.B2(n_400),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_546),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_485),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_510),
.B(n_514),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_542),
.B(n_519),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_508),
.C(n_503),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_549),
.B(n_553),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_499),
.C(n_501),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_536),
.C(n_534),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_555),
.B(n_563),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_558),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_541),
.C(n_545),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_498),
.C(n_488),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_523),
.B(n_504),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_567),
.B(n_568),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_531),
.C(n_524),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_574),
.B(n_585),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_551),
.B(n_535),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_577),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_555),
.B(n_537),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_578),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_519),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_579),
.B(n_584),
.Y(n_600)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_561),
.Y(n_580)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_580),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_581),
.B(n_548),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_570),
.Y(n_582)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_582),
.Y(n_599)
);

AOI322xp5_ASAP7_75t_L g583 ( 
.A1(n_562),
.A2(n_558),
.A3(n_565),
.B1(n_560),
.B2(n_520),
.C1(n_521),
.C2(n_571),
.Y(n_583)
);

BUFx24_ASAP7_75t_SL g606 ( 
.A(n_583),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_549),
.B(n_539),
.C(n_530),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_540),
.C(n_544),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_589),
.C(n_570),
.Y(n_601)
);

NAND5xp2_ASAP7_75t_L g587 ( 
.A(n_550),
.B(n_522),
.C(n_538),
.D(n_506),
.E(n_505),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_587),
.A2(n_554),
.B1(n_557),
.B2(n_564),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_567),
.B(n_381),
.C(n_389),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_560),
.A2(n_319),
.B1(n_354),
.B2(n_336),
.Y(n_590)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_590),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_576),
.B(n_569),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_591),
.B(n_593),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_573),
.B(n_556),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_596),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_587),
.A2(n_566),
.B1(n_550),
.B2(n_563),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_597),
.A2(n_607),
.B1(n_344),
.B2(n_395),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_601),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_584),
.B(n_568),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_605),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_572),
.A2(n_553),
.B(n_396),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_581),
.A2(n_586),
.B1(n_589),
.B2(n_582),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_592),
.B(n_575),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_609),
.B(n_610),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_579),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_588),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_611),
.B(n_619),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_607),
.B(n_601),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_613),
.B(n_617),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_597),
.A2(n_588),
.B1(n_336),
.B2(n_354),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_620),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_616),
.A2(n_344),
.B1(n_331),
.B2(n_314),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_606),
.A2(n_396),
.B(n_395),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_594),
.B(n_347),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_598),
.B(n_347),
.C(n_331),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_615),
.A2(n_595),
.B(n_599),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_622),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_594),
.C(n_596),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_603),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_630),
.C(n_624),
.Y(n_634)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_627),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_314),
.C(n_310),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_629),
.B(n_313),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_310),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_622),
.A2(n_618),
.B(n_612),
.Y(n_631)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_631),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_632),
.A2(n_636),
.B(n_637),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_634),
.A2(n_630),
.B1(n_628),
.B2(n_282),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_313),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_623),
.B(n_625),
.Y(n_637)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_638),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_635),
.A2(n_238),
.B(n_276),
.Y(n_639)
);

AOI31xp67_ASAP7_75t_SL g642 ( 
.A1(n_639),
.A2(n_276),
.A3(n_282),
.B(n_632),
.Y(n_642)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_642),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_641),
.C(n_643),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_646),
.B(n_640),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_633),
.Y(n_648)
);


endmodule