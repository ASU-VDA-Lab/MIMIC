module fake_jpeg_2362_n_489 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_489);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_489;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_7),
.B(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_61),
.Y(n_102)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_78),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_0),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_84),
.Y(n_142)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_48),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_24),
.B1(n_46),
.B2(n_45),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_98),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_99),
.A2(n_26),
.B(n_23),
.C(n_22),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_24),
.B1(n_46),
.B2(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_112),
.A2(n_120),
.B1(n_121),
.B2(n_131),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_135),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_27),
.B1(n_46),
.B2(n_45),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_57),
.B1(n_73),
.B2(n_53),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_67),
.B(n_27),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_35),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_72),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_139),
.B1(n_146),
.B2(n_153),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_75),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_70),
.B(n_48),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_37),
.C(n_36),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_26),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_42),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_25),
.C(n_31),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_77),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_32),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_154),
.B(n_26),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_105),
.A2(n_79),
.B1(n_76),
.B2(n_74),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g217 ( 
.A1(n_156),
.A2(n_159),
.B1(n_176),
.B2(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_160),
.Y(n_226)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_104),
.A2(n_69),
.B1(n_63),
.B2(n_56),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_162),
.Y(n_236)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_32),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_173),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_100),
.B(n_84),
.C(n_87),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_166),
.B(n_209),
.C(n_10),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_63),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_167),
.B(n_170),
.Y(n_219)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_56),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_177),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_32),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_112),
.A2(n_80),
.B1(n_25),
.B2(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_31),
.B1(n_58),
.B2(n_26),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_182),
.A2(n_210),
.B1(n_211),
.B2(n_119),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_122),
.Y(n_184)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_108),
.B(n_1),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_188),
.B(n_198),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_212),
.B1(n_133),
.B2(n_97),
.Y(n_230)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_191),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_99),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_195),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_1),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_98),
.B(n_99),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_199),
.B(n_206),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_121),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_124),
.B(n_119),
.Y(n_232)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_103),
.B(n_3),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g249 ( 
.A(n_207),
.B(n_208),
.Y(n_249)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_139),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_120),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_125),
.B(n_3),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_221),
.B(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_153),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_110),
.B1(n_130),
.B2(n_148),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_225),
.A2(n_231),
.B1(n_233),
.B2(n_240),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_253),
.B1(n_158),
.B2(n_164),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_110),
.B1(n_130),
.B2(n_148),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_SL g306 ( 
.A1(n_232),
.A2(n_249),
.B(n_216),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_125),
.B1(n_106),
.B2(n_138),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_138),
.A3(n_106),
.B1(n_97),
.B2(n_133),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_7),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_119),
.B1(n_9),
.B2(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_8),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_247),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_181),
.A2(n_8),
.B(n_9),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_243),
.A2(n_258),
.B(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_156),
.B(n_8),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_9),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_221),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_159),
.B(n_9),
.CI(n_10),
.CON(n_250),
.SN(n_250)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_250),
.B(n_263),
.C(n_215),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_254),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_176),
.B1(n_200),
.B2(n_207),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_167),
.B(n_10),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_256),
.C(n_170),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_13),
.C(n_14),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_211),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_263),
.B1(n_264),
.B2(n_217),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_174),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_208),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_192),
.A2(n_16),
.B1(n_17),
.B2(n_195),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_197),
.A2(n_17),
.B1(n_204),
.B2(n_170),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_295),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_184),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_272),
.C(n_277),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_218),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_228),
.A2(n_161),
.B1(n_201),
.B2(n_178),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_282),
.B1(n_283),
.B2(n_296),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_274),
.B(n_278),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_231),
.A2(n_169),
.B1(n_171),
.B2(n_185),
.Y(n_276)
);

OAI22x1_ASAP7_75t_L g346 ( 
.A1(n_276),
.A2(n_281),
.B1(n_296),
.B2(n_289),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_196),
.C(n_185),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_235),
.C(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_293),
.C(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_239),
.A2(n_247),
.B1(n_223),
.B2(n_245),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_217),
.B1(n_225),
.B2(n_219),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_292),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_244),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_305),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_224),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_290),
.B(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_241),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_261),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_214),
.B(n_233),
.C(n_216),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_217),
.A2(n_257),
.B1(n_264),
.B2(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_232),
.A2(n_250),
.B1(n_262),
.B2(n_226),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_299),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_250),
.A2(n_226),
.B1(n_258),
.B2(n_259),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_220),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_220),
.B(n_222),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_309),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_243),
.B(n_255),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_284),
.B(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_306),
.B(n_265),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_256),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_246),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_236),
.B(n_260),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_311),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_222),
.B(n_215),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_312),
.B(n_319),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_265),
.B1(n_244),
.B2(n_246),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_327),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_273),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_295),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_305),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_336),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_337),
.C(n_268),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_333),
.A2(n_348),
.B(n_284),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_334),
.B(n_349),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_246),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_293),
.C(n_270),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_275),
.B(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_345),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_344),
.B(n_266),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_275),
.B(n_282),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_299),
.B1(n_304),
.B2(n_303),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_283),
.B(n_307),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_297),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_269),
.B(n_272),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_279),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_352),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_320),
.B(n_269),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_353),
.B(n_364),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_357),
.A2(n_371),
.B(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_361),
.C(n_323),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_332),
.C(n_331),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_340),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_365),
.B1(n_368),
.B2(n_376),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_324),
.B(n_280),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_340),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_330),
.A2(n_347),
.B1(n_345),
.B2(n_325),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_373),
.B1(n_377),
.B2(n_371),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_277),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_336),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_291),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_381),
.Y(n_403)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_348),
.B(n_325),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_330),
.A2(n_281),
.B1(n_298),
.B2(n_309),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_377),
.A2(n_343),
.B1(n_342),
.B2(n_320),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_343),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_319),
.A2(n_322),
.B1(n_346),
.B2(n_327),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_338),
.B1(n_312),
.B2(n_334),
.Y(n_383)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_313),
.B1(n_338),
.B2(n_350),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_380),
.A2(n_355),
.B1(n_374),
.B2(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_382),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_383),
.A2(n_390),
.B1(n_394),
.B2(n_408),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_391),
.C(n_397),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_372),
.Y(n_388)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_338),
.B(n_329),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_389),
.A2(n_393),
.B(n_402),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_341),
.B1(n_313),
.B2(n_318),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_331),
.C(n_323),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_379),
.A2(n_343),
.B(n_328),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_318),
.B1(n_314),
.B2(n_315),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_360),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_404),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_315),
.C(n_342),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_372),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_356),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_378),
.C(n_375),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_407),
.C(n_365),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_363),
.B(n_375),
.C(n_371),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_409),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_403),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_414),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_398),
.B(n_362),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_413),
.B(n_415),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_408),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_393),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_374),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_368),
.C(n_380),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_427),
.C(n_428),
.Y(n_445)
);

XOR2x1_ASAP7_75t_SL g423 ( 
.A(n_401),
.B(n_380),
.Y(n_423)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_402),
.B(n_383),
.C(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_425),
.Y(n_434)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_380),
.C(n_358),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_SL g428 ( 
.A(n_407),
.B(n_355),
.C(n_359),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_399),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_431),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_370),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_416),
.A2(n_429),
.B1(n_411),
.B2(n_419),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_435),
.A2(n_418),
.B1(n_428),
.B2(n_425),
.Y(n_460)
);

OAI321xp33_ASAP7_75t_L g437 ( 
.A1(n_421),
.A2(n_430),
.A3(n_423),
.B1(n_424),
.B2(n_413),
.C(n_414),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_439),
.B1(n_446),
.B2(n_418),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_438),
.B(n_440),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_430),
.A2(n_390),
.B1(n_409),
.B2(n_394),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_386),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_444),
.B(n_447),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_389),
.B1(n_387),
.B2(n_385),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_443),
.A2(n_435),
.B1(n_447),
.B2(n_434),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_422),
.A2(n_387),
.B(n_385),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_420),
.A2(n_405),
.B1(n_381),
.B2(n_382),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_411),
.A2(n_404),
.B(n_376),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_395),
.Y(n_449)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_417),
.C(n_412),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_426),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_450),
.A2(n_455),
.B(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_452),
.A2(n_460),
.B1(n_437),
.B2(n_443),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_448),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_453),
.B(n_458),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_431),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_462),
.C(n_445),
.Y(n_469)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_448),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_433),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_412),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_461),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_427),
.C(n_391),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_471),
.C(n_454),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_453),
.A2(n_439),
.B1(n_433),
.B2(n_442),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_469),
.C(n_454),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_470),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_432),
.B1(n_445),
.B2(n_452),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_432),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_472),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_455),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_476),
.Y(n_482)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_474),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_451),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_466),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_480),
.B(n_481),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_477),
.C(n_478),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_484),
.A2(n_482),
.B1(n_463),
.B2(n_468),
.Y(n_485)
);

AOI321xp33_ASAP7_75t_L g486 ( 
.A1(n_485),
.A2(n_467),
.A3(n_463),
.B1(n_476),
.B2(n_459),
.C(n_483),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_SL g487 ( 
.A1(n_486),
.A2(n_467),
.B(n_460),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_462),
.B(n_450),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_457),
.Y(n_489)
);


endmodule