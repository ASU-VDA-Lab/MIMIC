module fake_jpeg_30525_n_516 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_72),
.Y(n_117)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_78),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_1),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_81),
.Y(n_145)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_3),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_101),
.Y(n_153)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_26),
.B(n_4),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_43),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_102),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_26),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_28),
.Y(n_138)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_46),
.B1(n_44),
.B2(n_53),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_118),
.A2(n_140),
.B1(n_161),
.B2(n_69),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_123),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_150),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_61),
.A2(n_46),
.B1(n_53),
.B2(n_36),
.Y(n_140)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_79),
.B(n_40),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_57),
.A2(n_23),
.B1(n_36),
.B2(n_53),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_72),
.B(n_40),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_164),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_171),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_117),
.A2(n_48),
.B(n_81),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_173),
.Y(n_264)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_176),
.Y(n_244)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_132),
.A2(n_53),
.B1(n_42),
.B2(n_23),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_137),
.B(n_104),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_146),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_198),
.Y(n_240)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_49),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_42),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_213),
.Y(n_229)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_43),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_117),
.A2(n_58),
.B1(n_103),
.B2(n_99),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_204),
.B1(n_221),
.B2(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_206),
.Y(n_252)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_202),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_125),
.A2(n_23),
.B1(n_51),
.B2(n_29),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_203),
.A2(n_205),
.B1(n_209),
.B2(n_212),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_75),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_169),
.B1(n_166),
.B2(n_51),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_52),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_208),
.Y(n_263)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_142),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_121),
.A2(n_66),
.B1(n_96),
.B2(n_94),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_210),
.A2(n_211),
.B1(n_77),
.B2(n_70),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_149),
.A2(n_65),
.B1(n_93),
.B2(n_92),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_140),
.A2(n_6),
.B(n_7),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_122),
.B(n_154),
.Y(n_226)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_39),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_223),
.Y(n_239)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_113),
.B(n_115),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_126),
.B1(n_109),
.B2(n_120),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_228),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_179),
.A2(n_138),
.B(n_112),
.C(n_29),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_227),
.B(n_255),
.Y(n_291)
);

OR2x2_ASAP7_75t_SL g228 ( 
.A(n_173),
.B(n_161),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_122),
.B1(n_148),
.B2(n_167),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_224),
.B1(n_209),
.B2(n_186),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_167),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_110),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_148),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_258),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_134),
.B1(n_126),
.B2(n_85),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_197),
.B1(n_188),
.B2(n_223),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_224),
.A2(n_47),
.B1(n_49),
.B2(n_45),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_47),
.B(n_52),
.C(n_39),
.Y(n_255)
);

NOR4xp25_ASAP7_75t_SL g257 ( 
.A(n_214),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_175),
.B(n_187),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_119),
.B1(n_151),
.B2(n_193),
.Y(n_267)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_119),
.B1(n_201),
.B2(n_222),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_269),
.A2(n_272),
.B1(n_236),
.B2(n_248),
.Y(n_319)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_228),
.B1(n_264),
.B2(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_278),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_206),
.B1(n_196),
.B2(n_171),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_280),
.Y(n_318)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_208),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_191),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_207),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_219),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_287),
.A2(n_295),
.B1(n_256),
.B2(n_238),
.Y(n_302)
);

AO22x1_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_240),
.B1(n_257),
.B2(n_249),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_218),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_212),
.B1(n_184),
.B2(n_183),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_294),
.B1(n_260),
.B2(n_237),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_240),
.A2(n_174),
.B1(n_220),
.B2(n_131),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_192),
.B1(n_172),
.B2(n_176),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_177),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_297),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_236),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_298),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_176),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_319),
.B1(n_311),
.B2(n_285),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_308),
.B1(n_316),
.B2(n_324),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_254),
.B(n_252),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_329),
.B(n_276),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_232),
.B1(n_253),
.B2(n_233),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_295),
.A2(n_244),
.B1(n_238),
.B2(n_243),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_309),
.A2(n_272),
.B1(n_287),
.B2(n_292),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_253),
.B(n_260),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_293),
.B(n_273),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_326),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_288),
.A2(n_245),
.B1(n_265),
.B2(n_235),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_263),
.B1(n_248),
.B2(n_261),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_227),
.C(n_234),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_268),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_255),
.B(n_243),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_334),
.B(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_275),
.Y(n_333)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_313),
.A2(n_266),
.B1(n_275),
.B2(n_276),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_337),
.B1(n_344),
.B2(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_313),
.A2(n_321),
.B1(n_301),
.B2(n_326),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_273),
.B(n_290),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_309),
.B(n_318),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_306),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_339),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_291),
.B(n_282),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_316),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_350),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_301),
.B1(n_325),
.B2(n_305),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_278),
.Y(n_345)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_302),
.B1(n_311),
.B2(n_294),
.Y(n_374)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_325),
.Y(n_365)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_284),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_279),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_353),
.A2(n_319),
.B1(n_318),
.B2(n_304),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_268),
.B(n_280),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_314),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_283),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_358),
.A2(n_359),
.B1(n_317),
.B2(n_323),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_320),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_339),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_362),
.A2(n_369),
.B1(n_371),
.B2(n_383),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_375),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_307),
.C(n_308),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_389),
.C(n_350),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_353),
.B1(n_318),
.B2(n_337),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_344),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_335),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_374),
.A2(n_246),
.B1(n_230),
.B2(n_202),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_323),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_333),
.B1(n_342),
.B2(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_343),
.A2(n_269),
.B1(n_267),
.B2(n_280),
.Y(n_383)
);

AOI21x1_ASAP7_75t_SL g384 ( 
.A1(n_354),
.A2(n_280),
.B(n_176),
.Y(n_384)
);

INVx13_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_332),
.A2(n_280),
.B(n_262),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_388),
.B(n_347),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_345),
.B(n_262),
.C(n_277),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_357),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_390),
.B(n_410),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_387),
.B(n_340),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_394),
.B(n_396),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_409),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_351),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_366),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_404),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_338),
.B(n_331),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_398),
.A2(n_379),
.B(n_360),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_352),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_399),
.A2(n_412),
.B(n_398),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_414),
.Y(n_417)
);

OAI32xp33_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_341),
.A3(n_358),
.B1(n_336),
.B2(n_330),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_359),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_406),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_375),
.C(n_378),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_346),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_368),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_377),
.B(n_33),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_413),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_389),
.B(n_270),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_234),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_415),
.A2(n_416),
.B1(n_381),
.B2(n_373),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_429),
.C(n_435),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_420),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_405),
.A2(n_363),
.B(n_388),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_399),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_374),
.B1(n_371),
.B2(n_369),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_426),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_401),
.B1(n_409),
.B2(n_402),
.Y(n_426)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_362),
.C(n_370),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_405),
.A2(n_383),
.B1(n_370),
.B2(n_380),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_401),
.B1(n_399),
.B2(n_403),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_380),
.C(n_386),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_408),
.B(n_376),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_408),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_441),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_395),
.C(n_391),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_445),
.C(n_450),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_400),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_404),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_423),
.A2(n_415),
.B(n_373),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_448),
.A2(n_421),
.B(n_433),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_416),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_411),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_430),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_419),
.C(n_434),
.Y(n_452)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_454),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_411),
.C(n_246),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_417),
.C(n_437),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_439),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_453),
.A2(n_431),
.B1(n_424),
.B2(n_426),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_472),
.Y(n_475)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_469),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_456),
.A2(n_420),
.B1(n_432),
.B2(n_422),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_468),
.Y(n_486)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_471),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_446),
.A2(n_417),
.B1(n_438),
.B2(n_427),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_455),
.A2(n_230),
.B1(n_45),
.B2(n_33),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_458),
.B(n_440),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_477),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_445),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_443),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_480),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_462),
.A2(n_440),
.B1(n_450),
.B2(n_444),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_482),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_28),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_8),
.B(n_9),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_108),
.C(n_9),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_470),
.C(n_10),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_472),
.Y(n_485)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_485),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_468),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_490),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_478),
.A2(n_486),
.B1(n_481),
.B2(n_469),
.Y(n_488)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_474),
.A2(n_467),
.B(n_463),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_492),
.B(n_486),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_484),
.A2(n_470),
.B(n_9),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_497),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_499),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_476),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_502),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_476),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_494),
.A2(n_8),
.B(n_11),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

AOI21xp33_ASAP7_75t_L g506 ( 
.A1(n_500),
.A2(n_491),
.B(n_488),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_498),
.B(n_503),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_510),
.C(n_508),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_495),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_507),
.B(n_490),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_11),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_12),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_13),
.C(n_14),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_13),
.C(n_14),
.Y(n_516)
);


endmodule