module real_aes_7683_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g188 ( .A1(n_0), .A2(n_189), .B(n_192), .C(n_196), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_1), .B(n_180), .Y(n_199) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g463 ( .A(n_2), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_3), .B(n_190), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_4), .A2(n_153), .B(n_156), .C(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_5), .A2(n_148), .B(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_6), .A2(n_148), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_7), .B(n_180), .Y(n_576) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_8), .A2(n_182), .B(n_254), .Y(n_253) );
AND2x6_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_10), .A2(n_153), .B(n_156), .C(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g537 ( .A(n_11), .Y(n_537) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_12), .B(n_39), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_13), .B(n_195), .Y(n_548) );
INVx1_ASAP7_75t_L g174 ( .A(n_14), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_15), .B(n_190), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_16), .A2(n_191), .B(n_556), .C(n_558), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_17), .B(n_180), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_18), .B(n_168), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_19), .A2(n_156), .B(n_159), .C(n_167), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_20), .A2(n_194), .B(n_262), .C(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_21), .B(n_195), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_22), .B(n_195), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_23), .Y(n_518) );
INVx1_ASAP7_75t_L g498 ( .A(n_24), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_25), .A2(n_156), .B(n_167), .C(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_26), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_27), .Y(n_544) );
INVx1_ASAP7_75t_L g512 ( .A(n_28), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_29), .A2(n_148), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g151 ( .A(n_30), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_31), .A2(n_206), .B(n_207), .C(n_211), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_32), .A2(n_33), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_32), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_33), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_34), .A2(n_194), .B(n_573), .C(n_575), .Y(n_572) );
INVxp67_ASAP7_75t_L g513 ( .A(n_35), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_36), .B(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_37), .A2(n_156), .B(n_167), .C(n_497), .Y(n_496) );
CKINVDCx14_ASAP7_75t_R g571 ( .A(n_38), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_40), .A2(n_196), .B(n_535), .C(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_41), .B(n_147), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_42), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_43), .B(n_190), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_44), .B(n_148), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_45), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_46), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_47), .A2(n_206), .B(n_211), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g193 ( .A(n_48), .Y(n_193) );
INVx1_ASAP7_75t_L g237 ( .A(n_49), .Y(n_237) );
INVx1_ASAP7_75t_L g584 ( .A(n_50), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_51), .B(n_148), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_52), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_53), .A2(n_105), .B1(n_117), .B2(n_772), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g533 ( .A(n_54), .Y(n_533) );
AOI22xp5_ASAP7_75t_SL g470 ( .A1(n_55), .A2(n_461), .B1(n_471), .B2(n_767), .Y(n_470) );
INVx1_ASAP7_75t_L g154 ( .A(n_56), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_57), .B(n_148), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_58), .B(n_180), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_59), .A2(n_166), .B(n_222), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g173 ( .A(n_60), .Y(n_173) );
INVx1_ASAP7_75t_SL g574 ( .A(n_61), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_62), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_63), .B(n_190), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_64), .B(n_180), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_65), .B(n_191), .Y(n_272) );
INVx1_ASAP7_75t_L g521 ( .A(n_66), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_67), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_68), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_69), .A2(n_156), .B(n_211), .C(n_220), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_70), .Y(n_246) );
INVx1_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_72), .A2(n_148), .B(n_532), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_73), .A2(n_95), .B1(n_133), .B2(n_134), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_73), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_74), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_75), .A2(n_103), .B1(n_480), .B2(n_481), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_75), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_76), .A2(n_148), .B(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_77), .A2(n_147), .B(n_508), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_78), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_79), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_79), .Y(n_477) );
INVx1_ASAP7_75t_L g554 ( .A(n_80), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_81), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_82), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_83), .A2(n_148), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g557 ( .A(n_84), .Y(n_557) );
INVx2_ASAP7_75t_L g171 ( .A(n_85), .Y(n_171) );
INVx1_ASAP7_75t_L g547 ( .A(n_86), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_87), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_88), .B(n_195), .Y(n_273) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
OR2x2_ASAP7_75t_L g460 ( .A(n_89), .B(n_461), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_90), .A2(n_156), .B(n_211), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_91), .B(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g208 ( .A(n_92), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_93), .B(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_L g249 ( .A(n_94), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_95), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_96), .A2(n_476), .B1(n_482), .B2(n_483), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_96), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_97), .B(n_182), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_98), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g221 ( .A(n_99), .Y(n_221) );
INVx1_ASAP7_75t_L g268 ( .A(n_100), .Y(n_268) );
INVx2_ASAP7_75t_L g587 ( .A(n_101), .Y(n_587) );
AND2x2_ASAP7_75t_L g239 ( .A(n_102), .B(n_170), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_103), .Y(n_480) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g772 ( .A(n_107), .Y(n_772) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g472 ( .A(n_113), .Y(n_472) );
INVx1_ASAP7_75t_L g485 ( .A(n_113), .Y(n_485) );
NOR2x2_ASAP7_75t_L g769 ( .A(n_113), .B(n_461), .Y(n_769) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_469), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g771 ( .A(n_122), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_458), .B(n_465), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_127), .B(n_181), .Y(n_549) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_135), .B2(n_136), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_135), .A2(n_136), .B1(n_474), .B2(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_413), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_348), .Y(n_137) );
NAND4xp25_ASAP7_75t_SL g138 ( .A(n_139), .B(n_293), .C(n_317), .D(n_340), .Y(n_138) );
AOI221xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_230), .B1(n_264), .B2(n_277), .C(n_280), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_200), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_142), .A2(n_178), .B1(n_231), .B2(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_142), .B(n_201), .Y(n_351) );
AND2x2_ASAP7_75t_L g370 ( .A(n_142), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_142), .B(n_354), .Y(n_440) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_178), .Y(n_142) );
AND2x2_ASAP7_75t_L g308 ( .A(n_143), .B(n_201), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_143), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g331 ( .A(n_143), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g336 ( .A(n_143), .B(n_179), .Y(n_336) );
INVx2_ASAP7_75t_L g368 ( .A(n_143), .Y(n_368) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_143), .Y(n_412) );
AND2x2_ASAP7_75t_L g429 ( .A(n_143), .B(n_306), .Y(n_429) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g347 ( .A(n_144), .B(n_306), .Y(n_347) );
AND2x4_ASAP7_75t_L g361 ( .A(n_144), .B(n_178), .Y(n_361) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_144), .Y(n_365) );
AND2x2_ASAP7_75t_L g385 ( .A(n_144), .B(n_300), .Y(n_385) );
AND2x2_ASAP7_75t_L g435 ( .A(n_144), .B(n_202), .Y(n_435) );
AND2x2_ASAP7_75t_L g445 ( .A(n_144), .B(n_179), .Y(n_445) );
OR2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_175), .Y(n_144) );
AOI21xp5_ASAP7_75t_SL g145 ( .A1(n_146), .A2(n_155), .B(n_168), .Y(n_145) );
BUFx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_149), .B(n_153), .Y(n_269) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g263 ( .A(n_151), .Y(n_263) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx3_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx1_ASAP7_75t_L g259 ( .A(n_152), .Y(n_259) );
BUFx3_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
INVx4_ASAP7_75t_SL g198 ( .A(n_153), .Y(n_198) );
INVx5_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_157), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_165), .Y(n_159) );
INVx2_ASAP7_75t_L g164 ( .A(n_161), .Y(n_164) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_208), .B(n_209), .C(n_210), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_210), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_164), .A2(n_521), .B(n_522), .C(n_523), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_164), .A2(n_523), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_165), .A2(n_190), .B(n_498), .C(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_166), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_169), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g177 ( .A(n_170), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_170), .A2(n_234), .B(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_170), .A2(n_269), .B(n_495), .C(n_496), .Y(n_494) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_170), .A2(n_531), .B(n_538), .Y(n_530) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_171), .B(n_172), .Y(n_170) );
AND2x2_ASAP7_75t_L g183 ( .A(n_171), .B(n_172), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_177), .A2(n_543), .B(n_549), .Y(n_542) );
AND2x2_ASAP7_75t_L g301 ( .A(n_178), .B(n_201), .Y(n_301) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_178), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_178), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g391 ( .A(n_178), .Y(n_391) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g279 ( .A(n_179), .B(n_216), .Y(n_279) );
AND2x2_ASAP7_75t_L g306 ( .A(n_179), .B(n_217), .Y(n_306) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_184), .B(n_199), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_181), .B(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_181), .A2(n_218), .B(n_228), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_181), .B(n_229), .Y(n_228) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_181), .A2(n_267), .B(n_274), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_181), .B(n_501), .Y(n_500) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_181), .A2(n_517), .B(n_524), .Y(n_516) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_182), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_182), .A2(n_255), .B(n_256), .Y(n_254) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_198), .Y(n_185) );
INVx2_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_187), .A2(n_198), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_187), .A2(n_198), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_187), .A2(n_198), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_187), .A2(n_198), .B(n_554), .C(n_555), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_187), .A2(n_198), .B(n_571), .C(n_572), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_SL g583 ( .A1(n_187), .A2(n_198), .B(n_584), .C(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g511 ( .A1(n_190), .A2(n_223), .B1(n_512), .B2(n_513), .Y(n_511) );
INVx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_191), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_194), .B(n_574), .Y(n_573) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g535 ( .A(n_195), .Y(n_535) );
INVx2_ASAP7_75t_L g523 ( .A(n_196), .Y(n_523) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_197), .Y(n_210) );
INVx1_ASAP7_75t_L g558 ( .A(n_197), .Y(n_558) );
INVx1_ASAP7_75t_L g211 ( .A(n_198), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_200), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_214), .Y(n_200) );
OR2x2_ASAP7_75t_L g332 ( .A(n_201), .B(n_215), .Y(n_332) );
AND2x2_ASAP7_75t_L g369 ( .A(n_201), .B(n_279), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_201), .B(n_300), .Y(n_380) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_201), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_201), .B(n_336), .Y(n_453) );
INVx5_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g278 ( .A(n_202), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_202), .B(n_215), .Y(n_287) );
AND2x2_ASAP7_75t_L g403 ( .A(n_202), .B(n_298), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_202), .B(n_336), .Y(n_425) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_212), .Y(n_202) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_215), .Y(n_371) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_216), .Y(n_323) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g300 ( .A(n_217), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_224), .C(n_225), .Y(n_220) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_223), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_223), .B(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g575 ( .A(n_226), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_240), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_231), .B(n_313), .Y(n_432) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_232), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g284 ( .A(n_232), .B(n_285), .Y(n_284) );
INVx5_ASAP7_75t_SL g292 ( .A(n_232), .Y(n_292) );
OR2x2_ASAP7_75t_L g315 ( .A(n_232), .B(n_285), .Y(n_315) );
OR2x2_ASAP7_75t_L g325 ( .A(n_232), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g388 ( .A(n_232), .B(n_242), .Y(n_388) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_232), .B(n_241), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g447 ( .A(n_232), .B(n_368), .C(n_448), .D(n_449), .Y(n_447) );
AND2x2_ASAP7_75t_L g457 ( .A(n_232), .B(n_289), .Y(n_457) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g282 ( .A(n_241), .B(n_278), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_241), .B(n_284), .Y(n_451) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
OR2x2_ASAP7_75t_L g291 ( .A(n_242), .B(n_292), .Y(n_291) );
INVx3_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_242), .B(n_266), .Y(n_310) );
INVxp67_ASAP7_75t_L g313 ( .A(n_242), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_242), .B(n_285), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_242), .B(n_252), .Y(n_379) );
AND2x2_ASAP7_75t_L g394 ( .A(n_242), .B(n_289), .Y(n_394) );
OR2x2_ASAP7_75t_L g423 ( .A(n_242), .B(n_252), .Y(n_423) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_250), .Y(n_242) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_243), .A2(n_552), .B(n_559), .Y(n_551) );
OA21x2_ASAP7_75t_L g568 ( .A1(n_243), .A2(n_569), .B(n_576), .Y(n_568) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_243), .A2(n_582), .B(n_588), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_251), .B(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_251), .B(n_292), .Y(n_431) );
OR2x2_ASAP7_75t_L g452 ( .A(n_251), .B(n_329), .Y(n_452) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g265 ( .A(n_252), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g289 ( .A(n_252), .B(n_285), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_252), .B(n_266), .Y(n_304) );
AND2x2_ASAP7_75t_L g374 ( .A(n_252), .B(n_298), .Y(n_374) );
AND2x2_ASAP7_75t_L g408 ( .A(n_252), .B(n_292), .Y(n_408) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_253), .B(n_292), .Y(n_311) );
AND2x2_ASAP7_75t_L g339 ( .A(n_253), .B(n_266), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_261), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_261), .A2(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_264), .B(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_265), .A2(n_354), .B1(n_390), .B2(n_407), .C(n_409), .Y(n_406) );
INVx5_ASAP7_75t_SL g285 ( .A(n_266), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_270), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_269), .A2(n_518), .B(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_269), .A2(n_544), .B(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g506 ( .A(n_276), .Y(n_506) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OAI33xp33_ASAP7_75t_L g305 ( .A1(n_278), .A2(n_306), .A3(n_307), .B1(n_309), .B2(n_312), .B3(n_316), .Y(n_305) );
OR2x2_ASAP7_75t_L g321 ( .A(n_278), .B(n_322), .Y(n_321) );
AOI322xp5_ASAP7_75t_L g430 ( .A1(n_278), .A2(n_347), .A3(n_354), .B1(n_431), .B2(n_432), .C1(n_433), .C2(n_436), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_278), .B(n_306), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_SL g454 ( .A1(n_278), .A2(n_306), .B(n_455), .C(n_457), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_279), .A2(n_294), .B1(n_299), .B2(n_302), .C(n_305), .Y(n_293) );
INVx1_ASAP7_75t_L g386 ( .A(n_279), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_279), .B(n_435), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B1(n_286), .B2(n_288), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g363 ( .A(n_284), .B(n_298), .Y(n_363) );
AND2x2_ASAP7_75t_L g421 ( .A(n_284), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g329 ( .A(n_285), .B(n_292), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_285), .B(n_298), .Y(n_357) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_287), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_287), .B(n_365), .Y(n_419) );
OAI321xp33_ASAP7_75t_L g438 ( .A1(n_287), .A2(n_360), .A3(n_439), .B1(n_440), .B2(n_441), .C(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g405 ( .A(n_288), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_289), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g344 ( .A(n_289), .B(n_292), .Y(n_344) );
AOI321xp33_ASAP7_75t_L g402 ( .A1(n_289), .A2(n_306), .A3(n_403), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_304), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_292), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_292), .B(n_378), .Y(n_415) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g338 ( .A(n_296), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g303 ( .A(n_297), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_301), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g334 ( .A(n_306), .Y(n_334) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_308), .B(n_343), .Y(n_392) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
OR2x2_ASAP7_75t_L g356 ( .A(n_311), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g401 ( .A(n_311), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_312), .A2(n_359), .B1(n_362), .B2(n_364), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g456 ( .A(n_315), .B(n_379), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_324), .B2(n_330), .C(n_333), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_SL g400 ( .A(n_326), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_328), .B(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_328), .A2(n_396), .B(n_398), .Y(n_395) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g441 ( .A(n_329), .B(n_423), .Y(n_441) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g343 ( .A(n_332), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g387 ( .A(n_339), .B(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g449 ( .A(n_339), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B(n_345), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_343), .B(n_361), .Y(n_397) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
NAND5xp2_ASAP7_75t_L g348 ( .A(n_349), .B(n_366), .C(n_375), .D(n_395), .E(n_402), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B(n_355), .C(n_358), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g390 ( .A(n_354), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_362), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
OAI21xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_370), .B(n_372), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_367), .A2(n_421), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_420) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AOI321xp33_ASAP7_75t_L g375 ( .A1(n_368), .A2(n_376), .A3(n_380), .B1(n_381), .B2(n_387), .C(n_389), .Y(n_375) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g446 ( .A(n_380), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g398 ( .A(n_383), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NOR2xp67_ASAP7_75t_SL g410 ( .A(n_384), .B(n_391), .Y(n_410) );
AOI321xp33_ASAP7_75t_SL g442 ( .A1(n_387), .A2(n_443), .A3(n_444), .B1(n_445), .B2(n_446), .C(n_447), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_392), .C(n_393), .Y(n_389) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_400), .B(n_408), .Y(n_437) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_412), .Y(n_409) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_438), .C(n_450), .Y(n_413) );
OAI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_420), .C(n_430), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_419), .A2(n_451), .B1(n_452), .B2(n_453), .C(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g443 ( .A(n_441), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g468 ( .A(n_460), .Y(n_468) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_465), .A2(n_470), .B(n_770), .Y(n_469) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_484), .B2(n_486), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_474), .A2(n_475), .B1(n_487), .B2(n_488), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g483 ( .A(n_476), .Y(n_483) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR4x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_657), .C(n_704), .D(n_744), .Y(n_488) );
NAND3xp33_ASAP7_75t_SL g489 ( .A(n_490), .B(n_603), .C(n_632), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_526), .B(n_560), .C(n_596), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_491), .A2(n_616), .B(n_633), .C(n_637), .Y(n_632) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_493), .B(n_595), .Y(n_594) );
INVx3_ASAP7_75t_SL g599 ( .A(n_493), .Y(n_599) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_493), .Y(n_611) );
AND2x4_ASAP7_75t_L g615 ( .A(n_493), .B(n_567), .Y(n_615) );
AND2x2_ASAP7_75t_L g626 ( .A(n_493), .B(n_516), .Y(n_626) );
OR2x2_ASAP7_75t_L g650 ( .A(n_493), .B(n_563), .Y(n_650) );
AND2x2_ASAP7_75t_L g663 ( .A(n_493), .B(n_568), .Y(n_663) );
AND2x2_ASAP7_75t_L g703 ( .A(n_493), .B(n_689), .Y(n_703) );
AND2x2_ASAP7_75t_L g710 ( .A(n_493), .B(n_673), .Y(n_710) );
AND2x2_ASAP7_75t_L g740 ( .A(n_493), .B(n_503), .Y(n_740) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_502), .B(n_667), .Y(n_679) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_515), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_503), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g617 ( .A(n_503), .B(n_515), .Y(n_617) );
BUFx3_ASAP7_75t_L g625 ( .A(n_503), .Y(n_625) );
OR2x2_ASAP7_75t_L g646 ( .A(n_503), .B(n_529), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_503), .B(n_667), .Y(n_757) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .B(n_514), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_505), .A2(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g564 ( .A(n_507), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_514), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g610 ( .A(n_515), .Y(n_610) );
AND2x2_ASAP7_75t_L g673 ( .A(n_515), .B(n_568), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_515), .A2(n_676), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_675) );
AND2x2_ASAP7_75t_L g689 ( .A(n_515), .B(n_563), .Y(n_689) );
AND2x2_ASAP7_75t_L g715 ( .A(n_515), .B(n_599), .Y(n_715) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g595 ( .A(n_516), .B(n_568), .Y(n_595) );
BUFx2_ASAP7_75t_L g729 ( .A(n_516), .Y(n_729) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI32xp33_ASAP7_75t_L g695 ( .A1(n_527), .A2(n_656), .A3(n_670), .B1(n_696), .B2(n_697), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
AND2x2_ASAP7_75t_L g636 ( .A(n_528), .B(n_580), .Y(n_636) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g618 ( .A(n_529), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_529), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g690 ( .A(n_529), .B(n_580), .Y(n_690) );
AND2x2_ASAP7_75t_L g701 ( .A(n_529), .B(n_593), .Y(n_701) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g602 ( .A(n_530), .B(n_581), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_530), .B(n_581), .Y(n_606) );
AND2x2_ASAP7_75t_L g641 ( .A(n_530), .B(n_592), .Y(n_641) );
AND2x2_ASAP7_75t_L g648 ( .A(n_530), .B(n_550), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_530), .A2(n_599), .B(n_610), .C(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g707 ( .A(n_530), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_530), .B(n_541), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_539), .B(n_590), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_539), .B(n_606), .Y(n_696) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_550), .Y(n_540) );
AND2x2_ASAP7_75t_L g593 ( .A(n_541), .B(n_551), .Y(n_593) );
OR2x2_ASAP7_75t_L g608 ( .A(n_541), .B(n_551), .Y(n_608) );
AND2x2_ASAP7_75t_L g631 ( .A(n_541), .B(n_592), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_541), .Y(n_635) );
AND2x2_ASAP7_75t_L g654 ( .A(n_541), .B(n_591), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_541), .A2(n_619), .B1(n_665), .B2(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_541), .B(n_707), .Y(n_731) );
AND2x2_ASAP7_75t_L g746 ( .A(n_541), .B(n_606), .Y(n_746) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g578 ( .A(n_542), .Y(n_578) );
AND2x2_ASAP7_75t_L g620 ( .A(n_542), .B(n_551), .Y(n_620) );
AND2x2_ASAP7_75t_L g622 ( .A(n_542), .B(n_580), .Y(n_622) );
AND3x2_ASAP7_75t_L g684 ( .A(n_542), .B(n_648), .C(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g719 ( .A(n_550), .B(n_591), .Y(n_719) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g580 ( .A(n_551), .B(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_551), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_551), .B(n_590), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_551), .B(n_631), .C(n_707), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_577), .B1(n_589), .B2(n_594), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_563), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g671 ( .A(n_563), .Y(n_671) );
OAI31xp33_ASAP7_75t_L g687 ( .A1(n_566), .A2(n_688), .A3(n_689), .B(n_690), .Y(n_687) );
AND2x2_ASAP7_75t_L g712 ( .A(n_566), .B(n_599), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_566), .B(n_625), .Y(n_758) );
AND2x2_ASAP7_75t_L g667 ( .A(n_567), .B(n_599), .Y(n_667) );
AND2x2_ASAP7_75t_L g728 ( .A(n_567), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g598 ( .A(n_568), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g656 ( .A(n_568), .Y(n_656) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g677 ( .A(n_578), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_579), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AOI221x1_ASAP7_75t_SL g644 ( .A1(n_580), .A2(n_645), .B1(n_647), .B2(n_649), .C(n_651), .Y(n_644) );
INVx2_ASAP7_75t_L g592 ( .A(n_581), .Y(n_592) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_581), .Y(n_686) );
INVx1_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_590), .B(n_607), .Y(n_699) );
INVx1_ASAP7_75t_SL g762 ( .A(n_590), .Y(n_762) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g680 ( .A(n_593), .B(n_606), .Y(n_680) );
INVx1_ASAP7_75t_L g748 ( .A(n_594), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_594), .B(n_677), .Y(n_761) );
INVx2_ASAP7_75t_SL g600 ( .A(n_595), .Y(n_600) );
AND2x2_ASAP7_75t_L g643 ( .A(n_595), .B(n_599), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_595), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_595), .B(n_670), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_600), .B(n_601), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_598), .B(n_670), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_598), .B(n_625), .Y(n_766) );
OR2x2_ASAP7_75t_L g638 ( .A(n_599), .B(n_617), .Y(n_638) );
AND2x2_ASAP7_75t_L g737 ( .A(n_599), .B(n_728), .Y(n_737) );
OAI22xp5_ASAP7_75t_SL g612 ( .A1(n_600), .A2(n_613), .B1(n_618), .B2(n_621), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_600), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g660 ( .A(n_602), .B(n_608), .Y(n_660) );
INVx1_ASAP7_75t_L g724 ( .A(n_602), .Y(n_724) );
AOI311xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_609), .A3(n_611), .B(n_612), .C(n_623), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_607), .A2(n_739), .B1(n_751), .B2(n_754), .C(n_756), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_607), .B(n_762), .Y(n_764) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g661 ( .A(n_609), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_610), .A2(n_652), .B(n_653), .C(n_655), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_SL g720 ( .A1(n_614), .A2(n_616), .B(n_721), .C(n_722), .Y(n_720) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_615), .B(n_689), .Y(n_755) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_618), .A2(n_638), .B1(n_639), .B2(n_642), .C(n_644), .Y(n_637) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g640 ( .A(n_620), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g723 ( .A(n_620), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_624), .A2(n_682), .B(n_683), .C(n_687), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_625), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_625), .B(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g647 ( .A(n_631), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_635), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g749 ( .A(n_638), .Y(n_749) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_641), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g676 ( .A(n_641), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g753 ( .A(n_641), .Y(n_753) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g694 ( .A(n_643), .B(n_670), .Y(n_694) );
INVx1_ASAP7_75t_SL g688 ( .A(n_650), .Y(n_688) );
INVx1_ASAP7_75t_L g665 ( .A(n_656), .Y(n_665) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_675), .C(n_691), .Y(n_657) );
AOI322xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .A3(n_662), .B1(n_664), .B2(n_668), .C1(n_672), .C2(n_674), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_659), .A2(n_712), .B(n_713), .C(n_720), .Y(n_711) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_662), .A2(n_683), .B1(n_714), .B2(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g672 ( .A(n_670), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g709 ( .A(n_670), .B(n_710), .Y(n_709) );
AOI32xp33_ASAP7_75t_L g760 ( .A1(n_670), .A2(n_761), .A3(n_762), .B1(n_763), .B2(n_765), .Y(n_760) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g682 ( .A(n_673), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_673), .A2(n_726), .B1(n_730), .B2(n_732), .C(n_735), .Y(n_725) );
AND2x2_ASAP7_75t_L g739 ( .A(n_673), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g742 ( .A(n_677), .B(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g752 ( .A(n_677), .B(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g743 ( .A(n_686), .B(n_707), .Y(n_743) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_695), .C(n_698), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_708), .B(n_711), .C(n_725), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_719), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g734 ( .A(n_731), .Y(n_734) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_741), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI211xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_747), .B(n_750), .C(n_760), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
endmodule