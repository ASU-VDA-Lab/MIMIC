module fake_jpeg_28214_n_22 (n_0, n_3, n_2, n_1, n_22);

input n_0;
input n_3;
input n_2;
input n_1;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_4;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g4 ( 
.A(n_1),
.Y(n_4)
);

INVx1_ASAP7_75t_L g5 ( 
.A(n_1),
.Y(n_5)
);

INVx3_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx8_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx4_ASAP7_75t_SL g8 ( 
.A(n_7),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_10),
.C(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_0),
.Y(n_9)
);

XNOR2xp5_ASAP7_75t_SL g12 ( 
.A(n_9),
.B(n_7),
.Y(n_12)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_9),
.A2(n_6),
.B1(n_5),
.B2(n_4),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_12),
.B1(n_6),
.B2(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_12),
.C(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_5),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_2),
.B(n_3),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_8),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_18),
.B(n_19),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_10),
.B(n_8),
.C(n_1),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_20),
.B(n_3),
.C(n_2),
.D(n_10),
.Y(n_22)
);


endmodule