module fake_jpeg_3404_n_491 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_491);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_59),
.Y(n_200)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_65),
.Y(n_178)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_17),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_80),
.A2(n_95),
.B(n_106),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_15),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_84),
.B(n_103),
.Y(n_133)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_14),
.B(n_13),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_98),
.Y(n_143)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_104),
.B(n_107),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g105 ( 
.A(n_38),
.B(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_37),
.B(n_12),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_113),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_50),
.B1(n_35),
.B2(n_30),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_53),
.B(n_13),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_13),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_115),
.B(n_63),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_36),
.B(n_11),
.CON(n_116),
.SN(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_0),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_118),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_31),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_120),
.Y(n_164)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_123),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_126),
.A2(n_163),
.B1(n_189),
.B2(n_199),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_50),
.B1(n_35),
.B2(n_30),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_130),
.A2(n_138),
.B1(n_176),
.B2(n_190),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_48),
.B1(n_46),
.B2(n_31),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_136),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_50),
.B1(n_35),
.B2(n_29),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_26),
.B1(n_23),
.B2(n_33),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_144),
.A2(n_167),
.B1(n_169),
.B2(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_45),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_175),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_48),
.B1(n_46),
.B2(n_33),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_81),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_106),
.A2(n_44),
.B1(n_35),
.B2(n_19),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_76),
.A2(n_42),
.B1(n_36),
.B2(n_35),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_0),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_165),
.B(n_173),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_55),
.A2(n_19),
.B1(n_27),
.B2(n_36),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_59),
.A2(n_42),
.B1(n_49),
.B2(n_3),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_0),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_98),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_65),
.A2(n_42),
.B1(n_49),
.B2(n_4),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_89),
.B(n_1),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_82),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_73),
.B(n_3),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_49),
.C(n_6),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_134),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_10),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_129),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_88),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_92),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_69),
.A2(n_94),
.B1(n_103),
.B2(n_101),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_93),
.B(n_10),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_56),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_195),
.A2(n_203),
.B1(n_132),
.B2(n_172),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_7),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_154),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_116),
.A2(n_8),
.B1(n_41),
.B2(n_51),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_195),
.B1(n_192),
.B2(n_143),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_117),
.A2(n_84),
.B1(n_34),
.B2(n_43),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_95),
.A2(n_84),
.B1(n_115),
.B2(n_81),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_151),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_205),
.B(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_207),
.B(n_213),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_162),
.B(n_133),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_238),
.Y(n_287)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_216),
.Y(n_314)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_226),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_164),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_232),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_142),
.B(n_152),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_228),
.Y(n_323)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_128),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_231),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_131),
.B(n_151),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g233 ( 
.A(n_143),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_264),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_189),
.A2(n_170),
.B1(n_197),
.B2(n_145),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_252),
.B1(n_255),
.B2(n_261),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_124),
.B(n_194),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_241),
.Y(n_285)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_191),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_135),
.A2(n_139),
.B1(n_147),
.B2(n_146),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_242),
.A2(n_249),
.B1(n_253),
.B2(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_161),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_244),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_139),
.B(n_152),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_142),
.B(n_140),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_121),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_259),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_137),
.B(n_140),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_251),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_141),
.B(n_185),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_254),
.Y(n_298)
);

NAND2x1p5_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_158),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_126),
.A2(n_177),
.B1(n_186),
.B2(n_121),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_146),
.A2(n_155),
.B1(n_147),
.B2(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_196),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_177),
.A2(n_187),
.B1(n_122),
.B2(n_149),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_155),
.A2(n_172),
.B1(n_122),
.B2(n_144),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_168),
.A2(n_200),
.B1(n_125),
.B2(n_181),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_258),
.A2(n_256),
.B1(n_228),
.B2(n_230),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_174),
.B(n_196),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_187),
.A2(n_149),
.B1(n_200),
.B2(n_174),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_266),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_153),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_148),
.A2(n_159),
.B(n_151),
.C(n_197),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_265),
.A2(n_214),
.B(n_213),
.C(n_206),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_201),
.B(n_153),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_267),
.B(n_268),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_148),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_129),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_269),
.B(n_271),
.Y(n_306)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_143),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_272),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_153),
.Y(n_272)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_233),
.B1(n_264),
.B2(n_263),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_255),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_210),
.B1(n_236),
.B2(n_252),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_309),
.B1(n_237),
.B2(n_240),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_249),
.A2(n_250),
.B1(n_210),
.B2(n_209),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_308),
.B1(n_311),
.B2(n_319),
.Y(n_325)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_301),
.A2(n_296),
.B(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_209),
.A2(n_225),
.B1(n_223),
.B2(n_251),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_234),
.A2(n_221),
.B1(n_265),
.B2(n_238),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_251),
.A2(n_263),
.B1(n_247),
.B2(n_260),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_273),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_315),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_219),
.B(n_245),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_245),
.B(n_228),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_321),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_222),
.B(n_248),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_211),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_323),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_261),
.A2(n_218),
.B1(n_216),
.B2(n_259),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g342 ( 
.A1(n_324),
.A2(n_283),
.B(n_318),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_332),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_217),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_336),
.C(n_302),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_277),
.A2(n_275),
.B1(n_271),
.B2(n_231),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_330),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_309),
.A2(n_301),
.B(n_291),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_329),
.A2(n_335),
.B(n_350),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_274),
.B1(n_269),
.B2(n_208),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_331),
.A2(n_348),
.B1(n_357),
.B2(n_314),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_212),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_333),
.B(n_343),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_270),
.B(n_272),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_235),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_334),
.Y(n_368)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_299),
.B(n_320),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_344),
.B(n_352),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_276),
.A2(n_298),
.B1(n_292),
.B2(n_284),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_346),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_285),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_318),
.A2(n_320),
.B(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_276),
.A2(n_284),
.B(n_298),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_349),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_292),
.B1(n_313),
.B2(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_286),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_282),
.B(n_293),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_351),
.A2(n_356),
.B(n_280),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_304),
.B(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_279),
.B(n_303),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_359),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g356 ( 
.A1(n_282),
.A2(n_279),
.A3(n_303),
.B1(n_312),
.B2(n_280),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_302),
.A2(n_306),
.B1(n_324),
.B2(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_289),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_390),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_354),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_371),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_342),
.A2(n_300),
.B(n_297),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

AOI221xp5_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_337),
.B1(n_355),
.B2(n_339),
.C(n_345),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_336),
.B(n_310),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_370),
.C(n_388),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_310),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_295),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_381),
.B(n_387),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_343),
.Y(n_381)
);

AO21x1_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_340),
.B(n_332),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_352),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_344),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_300),
.B(n_297),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_295),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_305),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_389),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_289),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_412),
.Y(n_416)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_396),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_376),
.A2(n_325),
.B1(n_348),
.B2(n_338),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_376),
.B1(n_371),
.B2(n_364),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_341),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_400),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_355),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_361),
.B(n_374),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_375),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_403),
.Y(n_425)
);

OA21x2_ASAP7_75t_SL g434 ( 
.A1(n_404),
.A2(n_405),
.B(n_410),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_383),
.B(n_381),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_325),
.B1(n_338),
.B2(n_330),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_281),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_413),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_415),
.Y(n_437)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_407),
.A2(n_384),
.B(n_386),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_417),
.A2(n_431),
.B(n_433),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_390),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_421),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_370),
.C(n_382),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_422),
.C(n_429),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_382),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_361),
.C(n_388),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_426),
.A2(n_408),
.B(n_393),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_368),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_418),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_428),
.A2(n_432),
.B1(n_391),
.B2(n_379),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_362),
.C(n_364),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_407),
.A2(n_367),
.B(n_374),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_397),
.A2(n_391),
.B1(n_376),
.B2(n_398),
.Y(n_432)
);

BUFx12f_ASAP7_75t_SL g433 ( 
.A(n_402),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_437),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_438),
.B(n_444),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_450),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_441),
.A2(n_351),
.B1(n_430),
.B2(n_423),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_373),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_437),
.Y(n_445)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_445),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_362),
.C(n_365),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_449),
.C(n_451),
.Y(n_461)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_416),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_452),
.B1(n_427),
.B2(n_326),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_365),
.C(n_375),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_422),
.C(n_421),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_378),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_420),
.A2(n_408),
.B1(n_374),
.B2(n_379),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_453),
.A2(n_432),
.B1(n_428),
.B2(n_420),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_346),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_460),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_447),
.A2(n_351),
.B1(n_433),
.B2(n_417),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_459),
.A2(n_443),
.B(n_453),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_426),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_434),
.Y(n_462)
);

AOI21x1_ASAP7_75t_SL g467 ( 
.A1(n_462),
.A2(n_440),
.B(n_443),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_431),
.C(n_392),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_446),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_464),
.B(n_449),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_466),
.B(n_471),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_467),
.A2(n_457),
.B(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_472),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_469),
.A2(n_465),
.B(n_455),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_435),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_474),
.A2(n_455),
.B1(n_460),
.B2(n_351),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_476),
.A2(n_477),
.B(n_469),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_480),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_436),
.B1(n_328),
.B2(n_396),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_461),
.C(n_439),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_484),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_473),
.C(n_467),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_461),
.C(n_451),
.Y(n_484)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_486),
.A2(n_346),
.B(n_415),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_483),
.A2(n_475),
.B(n_474),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_478),
.C(n_442),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_488),
.A2(n_489),
.B1(n_485),
.B2(n_442),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_414),
.Y(n_491)
);


endmodule