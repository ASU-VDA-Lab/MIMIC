module fake_jpeg_29497_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_42),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_27),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_52),
.B1(n_48),
.B2(n_22),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx9p33_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_89),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_22),
.B1(n_53),
.B2(n_33),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_101),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_46),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_31),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_46),
.B1(n_47),
.B2(n_43),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_109),
.B1(n_62),
.B2(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_65),
.B1(n_68),
.B2(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_108),
.B1(n_119),
.B2(n_88),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_65),
.B1(n_68),
.B2(n_43),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_45),
.B1(n_50),
.B2(n_44),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_85),
.Y(n_113)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_62),
.B1(n_45),
.B2(n_50),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_124),
.Y(n_161)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_137),
.Y(n_149)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_135),
.B1(n_103),
.B2(n_109),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_47),
.B1(n_44),
.B2(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_108),
.B1(n_105),
.B2(n_118),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_79),
.B1(n_93),
.B2(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_142),
.Y(n_151)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_112),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_157),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_112),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_152),
.B(n_156),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_111),
.B(n_121),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_83),
.B1(n_97),
.B2(n_118),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_139),
.B1(n_133),
.B2(n_138),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_104),
.B(n_79),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_104),
.C(n_82),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_78),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_163),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_114),
.B(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_114),
.B(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_170),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_186),
.B1(n_153),
.B2(n_160),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_181),
.Y(n_188)
);

INVx6_ASAP7_75t_SL g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_180),
.Y(n_193)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_98),
.B(n_114),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_78),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_90),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_29),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_26),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_146),
.C(n_161),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_191),
.C(n_196),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_189),
.B(n_26),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_146),
.C(n_158),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_157),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_200),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_155),
.B1(n_148),
.B2(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_125),
.B1(n_107),
.B2(n_142),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_150),
.C(n_162),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_183),
.B1(n_182),
.B2(n_166),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_145),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_145),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_164),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_80),
.B(n_61),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_214),
.B1(n_221),
.B2(n_229),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_213),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_212),
.B(n_30),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_168),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_180),
.B1(n_179),
.B2(n_171),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_134),
.B1(n_125),
.B2(n_131),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_216),
.B1(n_222),
.B2(n_80),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_141),
.B1(n_128),
.B2(n_83),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_117),
.B1(n_82),
.B2(n_73),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_141),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_190),
.B(n_128),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_128),
.B(n_73),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_226),
.B(n_86),
.Y(n_251)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_23),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_192),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_187),
.C(n_201),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_239),
.C(n_242),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_193),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_200),
.C(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_75),
.C(n_41),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_86),
.B(n_22),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_252),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_37),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_75),
.C(n_41),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_216),
.C(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_37),
.CI(n_30),
.CON(n_253),
.SN(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_61),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_86),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_218),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_258),
.B(n_264),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_221),
.B1(n_225),
.B2(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_224),
.C(n_225),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_274),
.C(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

BUFx12f_ASAP7_75t_SL g262 ( 
.A(n_236),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_266),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

BUFx12f_ASAP7_75t_SL g266 ( 
.A(n_253),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_270),
.B1(n_263),
.B2(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_245),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_244),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_28),
.C(n_35),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_234),
.C(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_284),
.C(n_273),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_246),
.C(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_40),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_289),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_240),
.B(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_3),
.B(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_72),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_272),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_72),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_5),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_300),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_256),
.C(n_258),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_275),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_302),
.B1(n_285),
.B2(n_304),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_268),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_35),
.B1(n_28),
.B2(n_49),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_33),
.B1(n_32),
.B2(n_9),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_4),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_35),
.C(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_276),
.B(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_279),
.C(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_316),
.C(n_302),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_314),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_5),
.C(n_6),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_72),
.C(n_30),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_323),
.Y(n_327)
);

OAI221xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_295),
.B1(n_8),
.B2(n_10),
.C(n_11),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_7),
.C(n_8),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_7),
.C(n_8),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_309),
.B(n_310),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_330),
.B1(n_322),
.B2(n_319),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_313),
.B(n_10),
.C(n_11),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_320),
.B(n_14),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_7),
.B(n_10),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_318),
.A3(n_32),
.B1(n_33),
.B2(n_14),
.C1(n_15),
.C2(n_12),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_327),
.C(n_14),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_12),
.C(n_32),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_32),
.B(n_33),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);


endmodule