module fake_jpeg_16919_n_388 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_47),
.B(n_59),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_53),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_15),
.B(n_14),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_0),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_34),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_79),
.B(n_104),
.Y(n_160)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_116),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_85),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_22),
.B1(n_20),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_84),
.A2(n_99),
.B1(n_17),
.B2(n_1),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_17),
.C(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_35),
.B1(n_29),
.B2(n_20),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_89),
.A2(n_96),
.B1(n_112),
.B2(n_124),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_35),
.B1(n_20),
.B2(n_40),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_35),
.B1(n_38),
.B2(n_19),
.Y(n_99)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_27),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_34),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_111),
.B(n_122),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_40),
.B1(n_41),
.B2(n_31),
.Y(n_112)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_40),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_41),
.B1(n_16),
.B2(n_21),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_51),
.B(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_37),
.B1(n_28),
.B2(n_32),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_78),
.B(n_19),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_47),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_132),
.B(n_8),
.Y(n_187)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_6),
.Y(n_179)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_91),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_141),
.Y(n_198)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_139),
.Y(n_218)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_41),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_142),
.B(n_146),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_31),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_32),
.B1(n_18),
.B2(n_31),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_159),
.B1(n_164),
.B2(n_167),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_152),
.Y(n_205)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_21),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_154),
.B(n_161),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_16),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_38),
.B1(n_17),
.B2(n_13),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_169),
.B1(n_9),
.B2(n_120),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_95),
.A2(n_12),
.B1(n_38),
.B2(n_2),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_170),
.B1(n_171),
.B2(n_138),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_171),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_112),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_1),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_177),
.Y(n_189)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_99),
.B1(n_133),
.B2(n_103),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_93),
.B(n_6),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_187),
.Y(n_229)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_84),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_191),
.A2(n_194),
.B1(n_209),
.B2(n_214),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_96),
.C(n_92),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_184),
.C(n_141),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_117),
.B(n_121),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_213),
.B(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_197),
.B(n_228),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_203),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_115),
.B(n_116),
.C(n_81),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_115),
.B1(n_117),
.B2(n_134),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_220),
.Y(n_244)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_123),
.B1(n_134),
.B2(n_81),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_143),
.A2(n_123),
.B1(n_119),
.B2(n_121),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_114),
.B1(n_119),
.B2(n_152),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_146),
.B(n_142),
.C(n_174),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_211),
.A2(n_190),
.B(n_230),
.C(n_210),
.Y(n_272)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_153),
.B(n_148),
.Y(n_213)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_162),
.B1(n_175),
.B2(n_157),
.Y(n_220)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_157),
.A2(n_185),
.B1(n_182),
.B2(n_158),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_222),
.B1(n_190),
.B2(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_168),
.A2(n_160),
.B1(n_172),
.B2(n_137),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_232),
.B1(n_207),
.B2(n_196),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_139),
.A2(n_136),
.B1(n_153),
.B2(n_150),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_239),
.C(n_255),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_186),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_240),
.B(n_242),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_186),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_253),
.C(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_247),
.B(n_251),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_230),
.B1(n_212),
.B2(n_201),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_226),
.C(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_192),
.CI(n_189),
.CON(n_255),
.SN(n_255)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_272),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_211),
.B(n_217),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_199),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_195),
.A2(n_202),
.B1(n_194),
.B2(n_220),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_252),
.B1(n_266),
.B2(n_243),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_204),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_193),
.B(n_201),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_208),
.B(n_198),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_191),
.A2(n_224),
.B(n_203),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_238),
.B(n_251),
.Y(n_298)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_200),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_200),
.B(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_293),
.B(n_297),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_230),
.B1(n_216),
.B2(n_233),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_281),
.B1(n_296),
.B2(n_248),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_233),
.B1(n_262),
.B2(n_244),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_239),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_282),
.B(n_292),
.Y(n_318)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_295),
.B1(n_283),
.B2(n_273),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_250),
.B(n_257),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_236),
.B1(n_249),
.B2(n_235),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_269),
.B(n_256),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_298),
.A2(n_278),
.B(n_301),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_240),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_237),
.Y(n_305)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_264),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_319),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_317),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_254),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_286),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_281),
.A2(n_264),
.B1(n_267),
.B2(n_258),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_270),
.B(n_258),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_288),
.B(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_320),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_283),
.A2(n_293),
.B1(n_291),
.B2(n_279),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_276),
.B(n_290),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_280),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_276),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_319),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_294),
.B(n_275),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_322),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_294),
.A2(n_275),
.B1(n_285),
.B2(n_277),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_300),
.B1(n_274),
.B2(n_286),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_295),
.B1(n_283),
.B2(n_149),
.Y(n_325)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_335),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_284),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_340),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_313),
.B1(n_310),
.B2(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_342),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_316),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_327),
.A2(n_310),
.B1(n_309),
.B2(n_307),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_344),
.A2(n_353),
.B1(n_355),
.B2(n_333),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_336),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_302),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_346),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_306),
.C(n_318),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_357),
.C(n_334),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_343),
.A2(n_312),
.B(n_321),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g366 ( 
.A1(n_354),
.A2(n_358),
.B(n_346),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_342),
.A2(n_318),
.B1(n_343),
.B2(n_330),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_341),
.C(n_338),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_337),
.B(n_341),
.Y(n_358)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_361),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_357),
.B(n_339),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_339),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_362),
.B(n_364),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_336),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_366),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_367),
.B(n_348),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_368),
.A2(n_349),
.B1(n_351),
.B2(n_353),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_373),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_360),
.C(n_364),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_375),
.B(n_376),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_371),
.B(n_351),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_370),
.Y(n_377)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

AOI322xp5_ASAP7_75t_L g381 ( 
.A1(n_378),
.A2(n_370),
.A3(n_374),
.B1(n_365),
.B2(n_349),
.C1(n_354),
.C2(n_346),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_382),
.B(n_379),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_384),
.A2(n_383),
.B(n_380),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_380),
.B(n_363),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_363),
.B(n_356),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_366),
.Y(n_388)
);


endmodule