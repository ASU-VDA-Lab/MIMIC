module fake_jpeg_1576_n_499 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_499);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_499;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_66),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_46),
.B1(n_36),
.B2(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_57),
.A2(n_26),
.B1(n_38),
.B2(n_33),
.Y(n_146)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_60),
.B(n_69),
.Y(n_145)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_14),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_75),
.Y(n_152)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_13),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_79),
.B(n_95),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_80),
.B(n_29),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_16),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_82),
.Y(n_139)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_86),
.B(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_10),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AND2x4_ASAP7_75t_SL g99 ( 
.A(n_29),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_29),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_43),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_107),
.B(n_131),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_36),
.B1(n_35),
.B2(n_24),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_108),
.A2(n_110),
.B1(n_19),
.B2(n_34),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_24),
.B1(n_35),
.B2(n_21),
.Y(n_110)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_41),
.B1(n_38),
.B2(n_26),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_88),
.B1(n_63),
.B2(n_76),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_29),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_77),
.A2(n_41),
.B1(n_44),
.B2(n_85),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_144),
.B1(n_78),
.B2(n_54),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_47),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_43),
.B1(n_33),
.B2(n_38),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_146),
.B1(n_20),
.B2(n_39),
.Y(n_183)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_49),
.Y(n_141)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_80),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_159),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_41),
.B1(n_29),
.B2(n_47),
.Y(n_144)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_51),
.B(n_42),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_161),
.B(n_154),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_162),
.B(n_158),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_172),
.Y(n_208)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_73),
.B1(n_65),
.B2(n_56),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_165),
.A2(n_183),
.B1(n_195),
.B2(n_157),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_26),
.B1(n_20),
.B2(n_50),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_186),
.B1(n_142),
.B2(n_123),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_167),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_78),
.C(n_54),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_196),
.C(n_206),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_177),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_105),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_175),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_20),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_188),
.Y(n_221)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_110),
.A2(n_50),
.B1(n_34),
.B2(n_19),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_0),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_1),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_199),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_34),
.C(n_19),
.Y(n_206)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_195),
.A2(n_112),
.B1(n_133),
.B2(n_108),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_217),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_125),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_214),
.B(n_228),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_120),
.C(n_134),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_112),
.B1(n_144),
.B2(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_230),
.B1(n_236),
.B2(n_240),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_235),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_168),
.A2(n_142),
.B1(n_147),
.B2(n_149),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_112),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_162),
.A2(n_119),
.B1(n_133),
.B2(n_151),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_189),
.A2(n_119),
.B1(n_126),
.B2(n_151),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_184),
.Y(n_251)
);

NAND2x1_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_129),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_196),
.B(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_242),
.B(n_221),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_173),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_196),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_165),
.B1(n_181),
.B2(n_185),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_248),
.A2(n_237),
.B1(n_210),
.B2(n_204),
.Y(n_302)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_254),
.Y(n_299)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_170),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_239),
.A2(n_179),
.B1(n_200),
.B2(n_197),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_260),
.B1(n_266),
.B2(n_269),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_175),
.B(n_187),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_261),
.B(n_232),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_263),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_194),
.B1(n_203),
.B2(n_201),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_193),
.B(n_198),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_212),
.A2(n_164),
.B(n_205),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_179),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_211),
.A2(n_182),
.B1(n_122),
.B2(n_101),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g268 ( 
.A(n_216),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_211),
.A2(n_116),
.B1(n_169),
.B2(n_171),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_171),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_270),
.B(n_225),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_218),
.A2(n_169),
.B1(n_190),
.B2(n_178),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_229),
.B1(n_215),
.B2(n_223),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_225),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_275),
.B(n_288),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_276),
.A2(n_281),
.B(n_282),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_217),
.C(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_254),
.C(n_247),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_243),
.B(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_286),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_232),
.B(n_213),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_230),
.B(n_211),
.C(n_219),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_283),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_246),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_243),
.A2(n_215),
.B1(n_223),
.B2(n_236),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_289),
.B1(n_300),
.B2(n_303),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_207),
.Y(n_288)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_253),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_290),
.Y(n_331)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_207),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_266),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_251),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_255),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_243),
.A2(n_242),
.B1(n_229),
.B2(n_210),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_272),
.B1(n_250),
.B2(n_256),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_243),
.A2(n_226),
.B1(n_222),
.B2(n_234),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_309),
.C(n_319),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_265),
.B1(n_250),
.B2(n_272),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_326),
.B1(n_279),
.B2(n_287),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_307),
.B(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_245),
.C(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_311),
.B(n_328),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_273),
.B(n_226),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_278),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_321),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_318),
.B(n_283),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_234),
.C(n_269),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_265),
.B1(n_259),
.B2(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_265),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_222),
.C(n_267),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_325),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_244),
.B1(n_249),
.B2(n_268),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_332),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_116),
.C(n_227),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_301),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_336),
.B(n_327),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_314),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_341),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_324),
.A2(n_314),
.B1(n_323),
.B2(n_333),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_343),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_313),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_313),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_362),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_333),
.B1(n_316),
.B2(n_325),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_284),
.B1(n_294),
.B2(n_304),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_358),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_306),
.A2(n_300),
.B1(n_303),
.B2(n_281),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_346),
.A2(n_348),
.B1(n_353),
.B2(n_360),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_305),
.B(n_291),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_309),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_326),
.B1(n_279),
.B2(n_276),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_304),
.A2(n_297),
.B1(n_282),
.B2(n_277),
.Y(n_358)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_319),
.A2(n_289),
.B1(n_282),
.B2(n_277),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_273),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_227),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_292),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_282),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_307),
.B(n_315),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_365),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_238),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_370),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_381),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_330),
.C(n_290),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_334),
.C(n_332),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_347),
.B(n_329),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_310),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_376),
.C(n_379),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_308),
.C(n_292),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_293),
.C(n_296),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_352),
.B(n_282),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_282),
.B(n_293),
.C(n_296),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_384),
.A2(n_358),
.B(n_354),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_238),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_386),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_249),
.C(n_252),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_268),
.B1(n_252),
.B2(n_257),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_389),
.B1(n_390),
.B2(n_380),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_233),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_391),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_339),
.A2(n_233),
.B(n_268),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_389),
.A2(n_390),
.B(n_346),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_257),
.B(n_121),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_121),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_371),
.A2(n_355),
.B1(n_360),
.B2(n_351),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_394),
.B1(n_409),
.B2(n_388),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_355),
.B1(n_351),
.B2(n_345),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_396),
.A2(n_405),
.B1(n_408),
.B2(n_410),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_403),
.B(n_387),
.Y(n_425)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_371),
.A2(n_357),
.B1(n_356),
.B2(n_354),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_413),
.B1(n_415),
.B2(n_391),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_357),
.B1(n_359),
.B2(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_349),
.B1(n_335),
.B2(n_113),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_386),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_378),
.A2(n_335),
.B1(n_113),
.B2(n_103),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_1),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_414),
.Y(n_434)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_1),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_378),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_376),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_417),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_373),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_375),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_423),
.Y(n_436)
);

INVx13_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_372),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_374),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_414),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_370),
.C(n_381),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_429),
.C(n_432),
.Y(n_447)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_382),
.C(n_366),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_176),
.B1(n_34),
.B2(n_3),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_430),
.A2(n_435),
.B1(n_394),
.B2(n_408),
.Y(n_437)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_407),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_431),
.B(n_1),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_1),
.C(n_2),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_399),
.B(n_396),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_412),
.B(n_400),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_404),
.A2(n_34),
.B1(n_2),
.B2(n_4),
.Y(n_435)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_427),
.A2(n_415),
.B1(n_401),
.B2(n_405),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_440),
.A2(n_442),
.B1(n_445),
.B2(n_448),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_425),
.A2(n_393),
.B1(n_399),
.B2(n_401),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_411),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_449),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_418),
.A2(n_413),
.B1(n_412),
.B2(n_403),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_438),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_410),
.B1(n_2),
.B2(n_4),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_423),
.C(n_416),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_426),
.C(n_424),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_453),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_421),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_420),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_457),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_429),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_463),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_450),
.B(n_432),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_461),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_2),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_9),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_464),
.B(n_466),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_5),
.C(n_6),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_446),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_9),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_447),
.B(n_5),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_438),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_440),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_477),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_436),
.C(n_439),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_478),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_455),
.A2(n_439),
.B(n_462),
.Y(n_474)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_474),
.A2(n_465),
.B(n_7),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_441),
.C(n_442),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_463),
.A2(n_443),
.B(n_6),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_SL g482 ( 
.A(n_479),
.B(n_459),
.C(n_460),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_457),
.C(n_468),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_483),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_482),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_476),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_487),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_475),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_471),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_475),
.B(n_9),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_486),
.C(n_470),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_478),
.C(n_469),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_491),
.A2(n_7),
.B(n_8),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_490),
.A2(n_485),
.B(n_481),
.Y(n_493)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_493),
.A2(n_494),
.B(n_495),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_492),
.B(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_7),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_8),
.B(n_497),
.Y(n_499)
);


endmodule