module fake_jpeg_27200_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_34),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_85)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_35),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_72),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_43),
.B1(n_44),
.B2(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_31),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_41),
.C(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_22),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_26),
.Y(n_100)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_89),
.Y(n_116)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_91),
.B1(n_44),
.B2(n_39),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_61),
.B1(n_48),
.B2(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_25),
.B1(n_22),
.B2(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_71),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_106),
.B1(n_109),
.B2(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_99),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_97),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_74),
.B1(n_84),
.B2(n_86),
.Y(n_120)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_18),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_39),
.B1(n_57),
.B2(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_126),
.B1(n_77),
.B2(n_80),
.Y(n_155)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_142),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_82),
.B1(n_84),
.B2(n_74),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_114),
.B1(n_108),
.B2(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_130),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_20),
.B(n_18),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_88),
.B1(n_63),
.B2(n_40),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_146),
.B1(n_70),
.B2(n_103),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_31),
.B1(n_34),
.B2(n_20),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_135),
.B(n_138),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_96),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_70),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_20),
.B(n_28),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_148),
.B(n_18),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_63),
.B1(n_40),
.B2(n_36),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_31),
.B(n_28),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_154),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_155),
.B1(n_172),
.B2(n_30),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_92),
.B(n_102),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_169),
.B(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_28),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_123),
.Y(n_183)
);

OA21x2_ASAP7_75t_R g154 ( 
.A1(n_122),
.A2(n_21),
.B(n_33),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_165),
.B1(n_168),
.B2(n_176),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_125),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_32),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_104),
.B1(n_103),
.B2(n_94),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_94),
.B1(n_36),
.B2(n_40),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_78),
.B(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_34),
.B1(n_29),
.B2(n_19),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_78),
.B1(n_29),
.B2(n_19),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_17),
.B1(n_19),
.B2(n_29),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_0),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_17),
.B1(n_21),
.B2(n_33),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_23),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_141),
.B(n_32),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_17),
.B1(n_21),
.B2(n_33),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_133),
.B(n_145),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_183),
.B(n_194),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_133),
.C(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_189),
.C(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_129),
.C(n_141),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_153),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_196),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_174),
.B1(n_150),
.B2(n_169),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_32),
.C(n_30),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_30),
.C(n_23),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_200),
.C(n_205),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_33),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_21),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_30),
.C(n_23),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_206),
.B1(n_179),
.B2(n_178),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_204),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_23),
.C(n_8),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_192),
.B1(n_212),
.B2(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_181),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_221),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_149),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_220),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_170),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_232),
.B1(n_201),
.B2(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_176),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_236),
.C(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_180),
.B(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_231),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_228),
.A2(n_191),
.B(n_159),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_230),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_196),
.B(n_165),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_210),
.B1(n_192),
.B2(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_172),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_159),
.C(n_168),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_237),
.B1(n_225),
.B2(n_215),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_258),
.B1(n_214),
.B2(n_226),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_187),
.B1(n_185),
.B2(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_252),
.Y(n_260)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_251),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_205),
.B1(n_200),
.B2(n_209),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_174),
.C(n_175),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_9),
.C(n_13),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_259),
.B(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_239),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_269),
.B1(n_274),
.B2(n_247),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_219),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_275),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_241),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_226),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_2),
.B(n_3),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_2),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_12),
.B(n_11),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_244),
.C(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_291),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_285),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_248),
.B1(n_242),
.B2(n_259),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_9),
.B1(n_10),
.B2(n_5),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_252),
.B(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_266),
.B1(n_268),
.B2(n_260),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_239),
.C(n_256),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_290),
.C(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_245),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_257),
.C(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_285),
.B1(n_286),
.B2(n_280),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_301),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_272),
.B(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_298),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_264),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_271),
.C(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_9),
.C(n_4),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_300),
.B(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_311),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_3),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_309),
.B(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_4),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_6),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_296),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_299),
.B(n_294),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_6),
.C(n_7),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_7),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_310),
.C(n_6),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_314),
.B(n_316),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_318),
.B(n_320),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_322),
.Y(n_328)
);


endmodule