module fake_jpeg_1818_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_23),
.B1(n_15),
.B2(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_23),
.B1(n_15),
.B2(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_45),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_32),
.B(n_23),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_31),
.B1(n_21),
.B2(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_22),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_8),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_37),
.C(n_10),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_70),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_35),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_69),
.C(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_5),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_48),
.Y(n_73)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_79),
.B(n_63),
.C(n_46),
.D(n_12),
.Y(n_87)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_72),
.B1(n_69),
.B2(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_79),
.B1(n_76),
.B2(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_81),
.B1(n_46),
.B2(n_12),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_88),
.B1(n_86),
.B2(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_85),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_0),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_89),
.C(n_91),
.Y(n_100)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_87),
.A3(n_12),
.B1(n_20),
.B2(n_24),
.C(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_1),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_20),
.B(n_1),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_99),
.C(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_2),
.Y(n_106)
);


endmodule