module fake_jpeg_20996_n_294 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_294);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_8),
.A2(n_2),
.B(n_9),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_27),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_49),
.C(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_21),
.B2(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_13),
.B(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_36),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_30),
.B(n_29),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_42),
.B(n_50),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_83),
.B1(n_84),
.B2(n_89),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_32),
.B1(n_34),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_34),
.B1(n_33),
.B2(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_39),
.B1(n_38),
.B2(n_41),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_46),
.B1(n_41),
.B2(n_33),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_47),
.C(n_30),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_46),
.B1(n_45),
.B2(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_85),
.B1(n_93),
.B2(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_112),
.Y(n_139)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_115),
.B(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_14),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_14),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OR2x6_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_74),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_96),
.C(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_126),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_108),
.B1(n_103),
.B2(n_110),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_75),
.B1(n_84),
.B2(n_96),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_84),
.B1(n_96),
.B2(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_137),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_96),
.B(n_1),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_135),
.B(n_138),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_89),
.B1(n_72),
.B2(n_52),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_16),
.B(n_28),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_0),
.C(n_1),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_1),
.C(n_2),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_99),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_109),
.B1(n_119),
.B2(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_127),
.B1(n_137),
.B2(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_107),
.B1(n_101),
.B2(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_155),
.B1(n_162),
.B2(n_165),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_151),
.B(n_158),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_152),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_113),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_115),
.B1(n_116),
.B2(n_112),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_164),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_113),
.B1(n_114),
.B2(n_106),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_163),
.B(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_142),
.B1(n_122),
.B2(n_132),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_114),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_131),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_139),
.B(n_26),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_108),
.B1(n_17),
.B2(n_25),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_123),
.B1(n_126),
.B2(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_180),
.B1(n_184),
.B2(n_158),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_174),
.A2(n_151),
.B(n_149),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_169),
.B1(n_146),
.B2(n_157),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_136),
.B1(n_120),
.B2(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_138),
.C(n_136),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_193),
.C(n_196),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_130),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_130),
.B1(n_135),
.B2(n_70),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_28),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_26),
.B1(n_17),
.B2(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_28),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_28),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_184),
.B1(n_172),
.B2(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_158),
.B(n_151),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_210),
.B(n_149),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_180),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_R g220 ( 
.A1(n_210),
.A2(n_179),
.B(n_178),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_227),
.CI(n_28),
.CON(n_240),
.SN(n_240)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_69),
.B1(n_68),
.B2(n_52),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_194),
.B(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_67),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_202),
.B(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_187),
.C(n_177),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.C(n_232),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_175),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_177),
.C(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_191),
.C(n_188),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_52),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_204),
.B1(n_211),
.B2(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_197),
.B1(n_192),
.B2(n_147),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_242),
.A3(n_243),
.B1(n_18),
.B2(n_223),
.C1(n_233),
.C2(n_6),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_147),
.C(n_173),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.C(n_67),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_2),
.B(n_3),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_245),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_218),
.Y(n_246)
);

OAI322xp33_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_219),
.A3(n_229),
.B1(n_231),
.B2(n_232),
.C1(n_226),
.C2(n_222),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_225),
.C(n_219),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_239),
.C(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_3),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_244),
.B(n_236),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_52),
.C(n_67),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_67),
.C(n_22),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_13),
.C(n_22),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_6),
.Y(n_273)
);

OAI211xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_255),
.B(n_7),
.C(n_9),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_243),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_22),
.B1(n_20),
.B2(n_8),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_255),
.B1(n_7),
.B2(n_8),
.Y(n_271)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_273),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_275),
.B1(n_276),
.B2(n_261),
.Y(n_280)
);

OR2x6_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_13),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_9),
.B(n_10),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_20),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_20),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_13),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_274),
.B1(n_260),
.B2(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_20),
.C(n_22),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_9),
.B(n_11),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.C(n_282),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_279),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_291),
.B(n_12),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_12),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_13),
.Y(n_294)
);


endmodule