module fake_jpeg_1731_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_40),
.C(n_53),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_41),
.C(n_47),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_44),
.B(n_42),
.C(n_46),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_48),
.B(n_2),
.C(n_3),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_49),
.B1(n_54),
.B2(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_73),
.B1(n_45),
.B2(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_43),
.B1(n_54),
.B2(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_61),
.B1(n_43),
.B2(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_41),
.B1(n_53),
.B2(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_84),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_62),
.C(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_86),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_48),
.C(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_50),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_0),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_73),
.Y(n_97)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_17),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_106),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_34),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_124),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_106),
.B(n_90),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_83),
.B1(n_80),
.B2(n_79),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_121),
.B1(n_122),
.B2(n_11),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_118),
.C(n_9),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_117),
.B1(n_12),
.B2(n_14),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_93),
.B1(n_99),
.B2(n_91),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_130),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_18),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_134),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_135),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_14),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_19),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_115),
.B(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_125),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_137),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_134),
.B(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_132),
.B1(n_128),
.B2(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_150),
.B(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_112),
.B1(n_129),
.B2(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_151),
.B(n_148),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_116),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_142),
.C(n_146),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_159),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_142),
.C(n_26),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_15),
.Y(n_162)
);


endmodule