module fake_jpeg_21313_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OR2x2_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_11),
.B1(n_15),
.B2(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_19),
.C(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_4),
.B(n_5),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_8),
.B(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_8),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.Y(n_40)
);

OAI221xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.C(n_30),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_39),
.C(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_21),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_21),
.Y(n_46)
);


endmodule