module real_aes_7818_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_83), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g438 ( .A(n_0), .Y(n_438) );
INVx1_ASAP7_75t_L g531 ( .A(n_1), .Y(n_531) );
INVx1_ASAP7_75t_L g148 ( .A(n_2), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_3), .A2(n_38), .B1(n_173), .B2(n_477), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g180 ( .A1(n_4), .A2(n_164), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_5), .B(n_162), .Y(n_543) );
AND2x6_ASAP7_75t_L g141 ( .A(n_6), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_8), .B(n_39), .Y(n_439) );
INVx1_ASAP7_75t_L g186 ( .A(n_9), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g133 ( .A(n_11), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_12), .B(n_154), .Y(n_486) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
INVx1_ASAP7_75t_L g525 ( .A(n_14), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_15), .B(n_129), .Y(n_514) );
AO32x2_ASAP7_75t_L g498 ( .A1(n_16), .A2(n_128), .A3(n_162), .B1(n_479), .B2(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_17), .B(n_173), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_18), .B(n_169), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_19), .B(n_129), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_20), .A2(n_49), .B1(n_173), .B2(n_477), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_21), .B(n_164), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_22), .A2(n_97), .B1(n_731), .B2(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_22), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_23), .A2(n_74), .B1(n_154), .B2(n_173), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_24), .B(n_173), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_25), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_26), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_28), .B(n_159), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_29), .B(n_152), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_30), .A2(n_86), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_30), .Y(n_119) );
INVx1_ASAP7_75t_L g201 ( .A(n_31), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_32), .B(n_159), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_33), .A2(n_444), .B1(n_729), .B2(n_730), .C1(n_733), .C2(n_735), .Y(n_443) );
INVx2_ASAP7_75t_L g139 ( .A(n_34), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_35), .B(n_173), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_36), .B(n_159), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_141), .B(n_144), .C(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g199 ( .A(n_40), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_41), .B(n_152), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_42), .B(n_173), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_43), .A2(n_84), .B1(n_221), .B2(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_44), .B(n_173), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_45), .B(n_173), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_46), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_47), .B(n_530), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_48), .B(n_164), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_50), .A2(n_59), .B1(n_154), .B2(n_173), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_51), .A2(n_144), .B1(n_154), .B2(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_52), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_53), .B(n_173), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_54), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_55), .B(n_173), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_56), .A2(n_172), .B(n_184), .C(n_185), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_57), .Y(n_234) );
INVx1_ASAP7_75t_L g182 ( .A(n_58), .Y(n_182) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_61), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_62), .B(n_173), .Y(n_532) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
AO32x2_ASAP7_75t_L g474 ( .A1(n_65), .A2(n_162), .A3(n_237), .B1(n_475), .B2(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g550 ( .A(n_66), .Y(n_550) );
INVx1_ASAP7_75t_L g465 ( .A(n_67), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_SL g168 ( .A1(n_68), .A2(n_169), .B(n_170), .C(n_172), .Y(n_168) );
INVxp67_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_70), .B(n_154), .Y(n_466) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_72), .Y(n_204) );
INVx1_ASAP7_75t_L g227 ( .A(n_73), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_75), .A2(n_141), .B(n_144), .C(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_76), .B(n_477), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_77), .B(n_154), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_78), .B(n_149), .Y(n_217) );
INVx2_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_80), .B(n_169), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_81), .B(n_154), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_82), .A2(n_141), .B(n_144), .C(n_147), .Y(n_143) );
OR2x2_ASAP7_75t_L g435 ( .A(n_83), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g447 ( .A(n_83), .B(n_437), .Y(n_447) );
INVx2_ASAP7_75t_L g452 ( .A(n_83), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_85), .A2(n_100), .B1(n_154), .B2(n_155), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_86), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_87), .B(n_159), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_88), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_89), .A2(n_141), .B(n_144), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_90), .Y(n_247) );
INVx1_ASAP7_75t_L g167 ( .A(n_91), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_92), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_93), .B(n_149), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_94), .A2(n_102), .B1(n_104), .B2(n_111), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_95), .B(n_154), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_96), .B(n_162), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_97), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_99), .A2(n_164), .B(n_165), .Y(n_163) );
BUFx4f_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_442), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g738 ( .A(n_113), .Y(n_738) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_433), .B(n_440), .Y(n_116) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g448 ( .A(n_121), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_121), .A2(n_449), .B1(n_454), .B2(n_734), .Y(n_733) );
NAND2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_349), .Y(n_121) );
NOR5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_272), .C(n_304), .D(n_319), .E(n_336), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_188), .B(n_209), .C(n_260), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_125), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_125), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_126), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_126), .B(n_206), .Y(n_273) );
AND2x2_ASAP7_75t_L g314 ( .A(n_126), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_126), .B(n_283), .Y(n_318) );
OR2x2_ASAP7_75t_L g355 ( .A(n_126), .B(n_194), .Y(n_355) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g193 ( .A(n_127), .B(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g263 ( .A(n_127), .Y(n_263) );
OR2x2_ASAP7_75t_L g426 ( .A(n_127), .B(n_266), .Y(n_426) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_156), .Y(n_127) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_128), .A2(n_195), .B(n_203), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_128), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g222 ( .A(n_128), .Y(n_222) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_130), .B(n_131), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_143), .Y(n_134) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_136), .A2(n_174), .B1(n_196), .B2(n_202), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_136), .A2(n_227), .B(n_228), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
AND2x4_ASAP7_75t_L g164 ( .A(n_137), .B(n_141), .Y(n_164) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g530 ( .A(n_138), .Y(n_530) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
INVx4_ASAP7_75t_SL g174 ( .A(n_141), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_141), .A2(n_464), .B(n_467), .Y(n_463) );
BUFx3_ASAP7_75t_L g479 ( .A(n_141), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_141), .A2(n_484), .B(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_141), .A2(n_524), .B(n_528), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_141), .A2(n_537), .B(n_540), .Y(n_536) );
INVx5_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
BUFx3_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
INVx1_ASAP7_75t_L g477 ( .A(n_145), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_151), .C(n_153), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_SL g464 ( .A1(n_149), .A2(n_172), .B(n_465), .C(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g501 ( .A(n_149), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_149), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_149), .A2(n_547), .B(n_548), .Y(n_546) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_150), .B(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_150), .B(n_186), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_150), .A2(n_152), .B1(n_476), .B2(n_478), .Y(n_475) );
INVx2_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx4_ASAP7_75t_L g243 ( .A(n_152), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_152), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_152), .A2(n_501), .B1(n_517), .B2(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_153), .A2(n_525), .B(n_526), .C(n_527), .Y(n_524) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_158), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_158), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g237 ( .A(n_159), .Y(n_237) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_159), .A2(n_463), .B(n_470), .Y(n_462) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_159), .A2(n_483), .B(n_491), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_160), .A2(n_329), .B1(n_330), .B2(n_333), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_160), .B(n_263), .Y(n_412) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_178), .Y(n_160) );
AND2x2_ASAP7_75t_L g208 ( .A(n_161), .B(n_194), .Y(n_208) );
AND2x2_ASAP7_75t_L g265 ( .A(n_161), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
INVx3_ASAP7_75t_L g283 ( .A(n_161), .Y(n_283) );
OR2x2_ASAP7_75t_L g303 ( .A(n_161), .B(n_266), .Y(n_303) );
AND2x2_ASAP7_75t_L g322 ( .A(n_161), .B(n_179), .Y(n_322) );
BUFx2_ASAP7_75t_L g354 ( .A(n_161), .Y(n_354) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_175), .Y(n_161) );
INVx4_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_162), .A2(n_536), .B(n_543), .Y(n_535) );
BUFx2_ASAP7_75t_L g251 ( .A(n_164), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_174), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_174), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_166), .A2(n_174), .B(n_253), .C(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g487 ( .A(n_169), .Y(n_487) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_176), .A2(n_180), .B(n_187), .Y(n_179) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_177), .B(n_224), .Y(n_223) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_177), .B(n_479), .C(n_516), .Y(n_515) );
AO21x1_ASAP7_75t_L g605 ( .A1(n_177), .A2(n_516), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g269 ( .A(n_178), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g192 ( .A(n_179), .Y(n_192) );
INVx2_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
OR2x2_ASAP7_75t_L g285 ( .A(n_179), .B(n_266), .Y(n_285) );
AND2x2_ASAP7_75t_L g315 ( .A(n_179), .B(n_194), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_179), .B(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g372 ( .A(n_179), .B(n_283), .Y(n_372) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_179), .B(n_208), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_184), .A2(n_489), .B(n_490), .Y(n_488) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_184), .A2(n_529), .B(n_550), .C(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp33_ASAP7_75t_SL g189 ( .A(n_190), .B(n_205), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_191), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_192), .A2(n_208), .B(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_192), .B(n_194), .Y(n_402) );
AND2x2_ASAP7_75t_L g338 ( .A(n_193), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_194), .Y(n_364) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g200 ( .A(n_198), .Y(n_200) );
INVx4_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_205), .B(n_263), .Y(n_431) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_206), .A2(n_374), .B1(n_375), .B2(n_380), .Y(n_373) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AND2x2_ASAP7_75t_L g264 ( .A(n_207), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g302 ( .A(n_207), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g339 ( .A(n_207), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_208), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g393 ( .A(n_208), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_235), .Y(n_210) );
INVx4_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
AND2x2_ASAP7_75t_L g357 ( .A(n_211), .B(n_324), .Y(n_357) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
INVx3_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
AND2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g294 ( .A(n_212), .Y(n_294) );
INVx2_ASAP7_75t_L g308 ( .A(n_212), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_212), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_212), .B(n_360), .Y(n_365) );
AND2x2_ASAP7_75t_L g430 ( .A(n_212), .B(n_400), .Y(n_430) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_219), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
INVx1_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_222), .A2(n_523), .B(n_533), .Y(n_522) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_222), .A2(n_545), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g271 ( .A(n_225), .B(n_249), .Y(n_271) );
INVx2_ASAP7_75t_L g291 ( .A(n_225), .Y(n_291) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_233), .Y(n_225) );
INVx1_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
AND2x2_ASAP7_75t_L g342 ( .A(n_235), .B(n_290), .Y(n_342) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
INVx2_ASAP7_75t_L g281 ( .A(n_236), .Y(n_281) );
INVx1_ASAP7_75t_L g289 ( .A(n_236), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_236), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_236), .B(n_291), .Y(n_345) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
AND2x2_ASAP7_75t_L g324 ( .A(n_248), .B(n_281), .Y(n_324) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
AND2x2_ASAP7_75t_L g360 ( .A(n_249), .B(n_291), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_255), .A2(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g527 ( .A(n_255), .Y(n_527) );
OAI21xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_267), .B(n_271), .Y(n_260) );
INVx1_ASAP7_75t_SL g305 ( .A(n_261), .Y(n_305) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_262), .B(n_269), .Y(n_362) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g311 ( .A(n_263), .B(n_266), .Y(n_311) );
AND2x2_ASAP7_75t_L g340 ( .A(n_263), .B(n_284), .Y(n_340) );
OR2x2_ASAP7_75t_L g343 ( .A(n_263), .B(n_303), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g407 ( .A1(n_264), .A2(n_356), .B1(n_408), .B2(n_409), .C1(n_411), .C2(n_413), .Y(n_407) );
BUFx2_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g310 ( .A(n_269), .B(n_311), .Y(n_310) );
INVx3_ASAP7_75t_SL g327 ( .A(n_269), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_269), .B(n_321), .Y(n_381) );
AND2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_276), .Y(n_316) );
INVx1_ASAP7_75t_L g335 ( .A(n_271), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_274), .B1(n_278), .B2(n_282), .C(n_286), .Y(n_272) );
OR2x2_ASAP7_75t_L g344 ( .A(n_274), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_299), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_276), .B(n_289), .Y(n_369) );
AND2x2_ASAP7_75t_L g374 ( .A(n_276), .B(n_324), .Y(n_374) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_276), .Y(n_384) );
NAND2x1_ASAP7_75t_SL g395 ( .A(n_276), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g280 ( .A(n_277), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_277), .B(n_295), .Y(n_326) );
INVx1_ASAP7_75t_L g392 ( .A(n_277), .Y(n_392) );
INVx1_ASAP7_75t_L g367 ( .A(n_278), .Y(n_367) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g379 ( .A(n_279), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_279), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g396 ( .A(n_280), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_280), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g299 ( .A(n_281), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_281), .B(n_291), .Y(n_312) );
INVx1_ASAP7_75t_L g378 ( .A(n_281), .Y(n_378) );
INVx1_ASAP7_75t_L g399 ( .A(n_282), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_292), .B(n_301), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x2_ASAP7_75t_L g432 ( .A(n_288), .B(n_365), .Y(n_432) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g400 ( .A(n_289), .B(n_360), .Y(n_400) );
AOI32xp33_ASAP7_75t_L g313 ( .A1(n_290), .A2(n_296), .A3(n_314), .B1(n_316), .B2(n_317), .Y(n_313) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_290), .A2(n_322), .A3(n_405), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g295 ( .A(n_291), .Y(n_295) );
INVx1_ASAP7_75t_L g405 ( .A(n_291), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_297), .B2(n_298), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_293), .B(n_299), .Y(n_348) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_294), .B(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g297 ( .A(n_295), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_295), .B(n_324), .Y(n_414) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_303), .B(n_398), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_306), .B1(n_309), .B2(n_312), .C(n_313), .Y(n_304) );
OR2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g359 ( .A(n_307), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g363 ( .A(n_317), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B1(n_325), .B2(n_327), .C(n_328), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_322), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_322), .Y(n_427) );
INVx1_ASAP7_75t_L g421 ( .A(n_324), .Y(n_421) );
INVx1_ASAP7_75t_SL g356 ( .A(n_325), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_327), .B(n_355), .Y(n_417) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g398 ( .A(n_332), .Y(n_398) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_341), .B1(n_343), .B2(n_344), .C(n_346), .Y(n_336) );
NOR2xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_338), .A2(n_356), .B1(n_402), .B2(n_403), .Y(n_401) );
CKINVDCx14_ASAP7_75t_R g341 ( .A(n_342), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_343), .A2(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR3xp33_ASAP7_75t_SL g349 ( .A(n_350), .B(n_382), .C(n_406), .Y(n_349) );
NAND4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_358), .C(n_366), .D(n_373), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
INVx3_ASAP7_75t_SL g423 ( .A(n_355), .Y(n_423) );
OR2x2_ASAP7_75t_L g428 ( .A(n_355), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_363), .B2(n_365), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_360), .B(n_378), .Y(n_419) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI21xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_370), .Y(n_366) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_388), .C(n_401), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g416 ( .A(n_387), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B1(n_394), .B2(n_397), .C1(n_399), .C2(n_400), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_SL g425 ( .A(n_398), .B(n_426), .C(n_427), .D(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_415), .C(n_424), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_424) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g441 ( .A(n_435), .Y(n_441) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_436), .B(n_452), .Y(n_737) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_440), .A2(n_443), .B(n_738), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_448), .B1(n_449), .B2(n_453), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g734 ( .A(n_446), .Y(n_734) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_650), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_599), .C(n_641), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_508), .B(n_553), .C(n_575), .Y(n_456) );
OAI211xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_471), .B(n_492), .C(n_503), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_459), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g662 ( .A(n_459), .B(n_579), .Y(n_662) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g564 ( .A(n_460), .B(n_495), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_460), .B(n_482), .Y(n_681) );
INVx1_ASAP7_75t_L g699 ( .A(n_460), .Y(n_699) );
AND2x2_ASAP7_75t_L g708 ( .A(n_460), .B(n_596), .Y(n_708) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g591 ( .A(n_461), .B(n_482), .Y(n_591) );
AND2x2_ASAP7_75t_L g649 ( .A(n_461), .B(n_596), .Y(n_649) );
INVx1_ASAP7_75t_L g693 ( .A(n_461), .Y(n_693) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g570 ( .A(n_462), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g578 ( .A(n_462), .Y(n_578) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_462), .Y(n_618) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .Y(n_472) );
AND2x2_ASAP7_75t_L g557 ( .A(n_473), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g590 ( .A(n_473), .Y(n_590) );
OR2x2_ASAP7_75t_L g716 ( .A(n_473), .B(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_473), .B(n_482), .Y(n_720) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
INVx1_ASAP7_75t_L g506 ( .A(n_474), .Y(n_506) );
AND2x2_ASAP7_75t_L g579 ( .A(n_474), .B(n_497), .Y(n_579) );
AND2x2_ASAP7_75t_L g619 ( .A(n_474), .B(n_498), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_479), .A2(n_546), .B(n_549), .Y(n_545) );
INVxp67_ASAP7_75t_L g661 ( .A(n_480), .Y(n_661) );
AND2x4_ASAP7_75t_L g686 ( .A(n_480), .B(n_579), .Y(n_686) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_481), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g496 ( .A(n_482), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g565 ( .A(n_482), .B(n_498), .Y(n_565) );
INVx1_ASAP7_75t_L g571 ( .A(n_482), .Y(n_571) );
INVx2_ASAP7_75t_L g597 ( .A(n_482), .Y(n_597) );
AND2x2_ASAP7_75t_L g613 ( .A(n_482), .B(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_493), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
AND2x2_ASAP7_75t_L g676 ( .A(n_495), .B(n_497), .Y(n_676) );
AND2x2_ASAP7_75t_L g593 ( .A(n_496), .B(n_578), .Y(n_593) );
AND2x2_ASAP7_75t_L g692 ( .A(n_496), .B(n_693), .Y(n_692) );
NOR2xp67_ASAP7_75t_L g614 ( .A(n_497), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g717 ( .A(n_497), .B(n_578), .Y(n_717) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g507 ( .A(n_498), .Y(n_507) );
AND2x2_ASAP7_75t_L g596 ( .A(n_498), .B(n_597), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_501), .A2(n_529), .B(n_531), .C(n_532), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_501), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g642 ( .A(n_505), .B(n_577), .Y(n_642) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_506), .B(n_578), .Y(n_627) );
INVx2_ASAP7_75t_L g626 ( .A(n_507), .Y(n_626) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_507), .A2(n_570), .B1(n_631), .B2(n_633), .C1(n_634), .C2(n_637), .Y(n_630) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g555 ( .A(n_512), .Y(n_555) );
OR2x2_ASAP7_75t_L g666 ( .A(n_512), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g588 ( .A(n_513), .Y(n_588) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_513), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g645 ( .A(n_513), .B(n_559), .Y(n_645) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g606 ( .A(n_514), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_519), .A2(n_609), .B1(n_648), .B2(n_649), .Y(n_647) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_534), .Y(n_519) );
INVx3_ASAP7_75t_L g581 ( .A(n_520), .Y(n_581) );
OR2x2_ASAP7_75t_L g714 ( .A(n_520), .B(n_590), .Y(n_714) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g587 ( .A(n_521), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g611 ( .A(n_521), .B(n_559), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_521), .B(n_535), .Y(n_667) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g558 ( .A(n_522), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g562 ( .A(n_522), .B(n_535), .Y(n_562) );
AND2x2_ASAP7_75t_L g638 ( .A(n_522), .B(n_585), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_522), .B(n_544), .Y(n_678) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_534), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g594 ( .A(n_534), .B(n_555), .Y(n_594) );
AND2x2_ASAP7_75t_L g598 ( .A(n_534), .B(n_588), .Y(n_598) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
INVx3_ASAP7_75t_L g559 ( .A(n_535), .Y(n_559) );
AND2x2_ASAP7_75t_L g584 ( .A(n_535), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g719 ( .A(n_535), .B(n_702), .Y(n_719) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_544), .Y(n_573) );
INVx2_ASAP7_75t_L g585 ( .A(n_544), .Y(n_585) );
AND2x2_ASAP7_75t_L g629 ( .A(n_544), .B(n_605), .Y(n_629) );
INVx1_ASAP7_75t_L g672 ( .A(n_544), .Y(n_672) );
OR2x2_ASAP7_75t_L g703 ( .A(n_544), .B(n_605), .Y(n_703) );
AND2x2_ASAP7_75t_L g723 ( .A(n_544), .B(n_559), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_556), .B(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g561 ( .A(n_555), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_555), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g680 ( .A(n_557), .Y(n_680) );
INVx2_ASAP7_75t_SL g574 ( .A(n_558), .Y(n_574) );
AND2x2_ASAP7_75t_L g694 ( .A(n_558), .B(n_588), .Y(n_694) );
INVx2_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_559), .B(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B1(n_566), .B2(n_572), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_562), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g728 ( .A(n_562), .Y(n_728) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g653 ( .A(n_564), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_564), .B(n_596), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_565), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g669 ( .A(n_565), .B(n_618), .Y(n_669) );
INVx2_ASAP7_75t_L g725 ( .A(n_565), .Y(n_725) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_568), .B(n_613), .Y(n_646) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_570), .B(n_590), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g707 ( .A(n_573), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_574), .A2(n_658), .B(n_660), .C(n_663), .Y(n_657) );
OR2x2_ASAP7_75t_L g684 ( .A(n_574), .B(n_588), .Y(n_684) );
OAI221xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_580), .B1(n_582), .B2(n_589), .C(n_592), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_577), .B(n_626), .Y(n_633) );
AND2x2_ASAP7_75t_L g675 ( .A(n_577), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g711 ( .A(n_577), .Y(n_711) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_578), .Y(n_602) );
INVx1_ASAP7_75t_L g615 ( .A(n_578), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g635 ( .A(n_581), .B(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g689 ( .A(n_581), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_581), .B(n_629), .Y(n_705) );
INVx2_ASAP7_75t_L g691 ( .A(n_582), .Y(n_691) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g632 ( .A(n_584), .B(n_603), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_584), .A2(n_600), .B(n_642), .C(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g610 ( .A(n_585), .B(n_605), .Y(n_610) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_589), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OR2x2_ASAP7_75t_L g658 ( .A(n_590), .B(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_598), .Y(n_592) );
INVx1_ASAP7_75t_L g712 ( .A(n_594), .Y(n_712) );
INVx1_ASAP7_75t_L g659 ( .A(n_596), .Y(n_659) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
AOI211xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_607), .C(n_630), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g622 ( .A(n_602), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g673 ( .A(n_603), .Y(n_673) );
AND2x2_ASAP7_75t_L g722 ( .A(n_603), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_612), .B(n_620), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g636 ( .A(n_610), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_610), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g628 ( .A(n_611), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g704 ( .A(n_611), .Y(n_704) );
OAI32xp33_ASAP7_75t_L g715 ( .A1(n_611), .A2(n_663), .A3(n_670), .B1(n_711), .B2(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_616), .Y(n_612) );
INVx1_ASAP7_75t_SL g683 ( .A(n_613), .Y(n_683) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g623 ( .A(n_619), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B(n_628), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_622), .A2(n_670), .B1(n_696), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_626), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g656 ( .A(n_640), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_647), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_649), .A2(n_691), .B1(n_692), .B2(n_694), .C(n_695), .Y(n_690) );
NAND5xp2_ASAP7_75t_L g650 ( .A(n_651), .B(n_674), .C(n_690), .D(n_700), .E(n_718), .Y(n_650) );
AOI211xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_654), .B(n_657), .C(n_664), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g721 ( .A(n_658), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_668), .B2(n_670), .Y(n_664) );
INVx1_ASAP7_75t_SL g697 ( .A(n_667), .Y(n_697) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_670), .A2(n_680), .A3(n_681), .B1(n_682), .B2(n_683), .C1(n_684), .C2(n_685), .Y(n_679) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g682 ( .A(n_672), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_672), .B(n_697), .Y(n_696) );
AOI211xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_677), .B(n_679), .C(n_687), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_683), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g726 ( .A(n_693), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_708), .B1(n_709), .B2(n_713), .C(n_715), .Y(n_700) );
OAI211xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_704), .B(n_705), .C(n_706), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g727 ( .A(n_703), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .C(n_724), .Y(n_718) );
AOI21xp33_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_726), .B(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
endmodule