module fake_jpeg_9598_n_31 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_29;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_10),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_5),
.B1(n_8),
.B2(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_0),
.B(n_2),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_24),
.C(n_14),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_21),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_19),
.B1(n_20),
.B2(n_13),
.Y(n_31)
);


endmodule