module real_jpeg_2637_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_58;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_51;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_71;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_70;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_5),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_17),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_8),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_52),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_32),
.B(n_51),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_25),
.B(n_31),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_18),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_62),
.Y(n_61)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_24),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_40),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_40),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_36),
.B(n_38),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_72),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_71),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_71),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);


endmodule