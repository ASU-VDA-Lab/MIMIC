module fake_aes_3924_n_951 (n_120, n_136, n_260, n_155, n_107, n_103, n_157, n_52, n_162, n_114, n_156, n_154, n_50, n_7, n_239, n_222, n_253, n_3, n_34, n_142, n_231, n_25, n_9, n_163, n_96, n_204, n_72, n_77, n_90, n_169, n_178, n_214, n_227, n_180, n_250, n_99, n_43, n_73, n_190, n_62, n_167, n_97, n_229, n_133, n_199, n_268, n_33, n_192, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_189, n_216, n_153, n_187, n_226, n_66, n_88, n_46, n_121, n_174, n_240, n_188, n_108, n_161, n_37, n_122, n_165, n_224, n_18, n_247, n_65, n_87, n_207, n_5, n_197, n_81, n_211, n_85, n_112, n_215, n_264, n_102, n_172, n_47, n_109, n_198, n_1, n_201, n_16, n_78, n_95, n_217, n_40, n_68, n_105, n_210, n_251, n_36, n_228, n_259, n_11, n_244, n_115, n_270, n_225, n_179, n_208, n_237, n_252, n_15, n_168, n_271, n_139, n_152, n_151, n_71, n_117, n_238, n_176, n_70, n_256, n_94, n_2, n_194, n_17, n_221, n_58, n_195, n_113, n_242, n_209, n_241, n_20, n_84, n_130, n_266, n_12, n_56, n_80, n_223, n_67, n_116, n_22, n_118, n_19, n_233, n_257, n_202, n_26, n_203, n_261, n_243, n_39, n_101, n_98, n_150, n_220, n_235, n_38, n_230, n_245, n_104, n_100, n_159, n_24, n_141, n_35, n_91, n_146, n_160, n_32, n_148, n_149, n_246, n_263, n_93, n_191, n_143, n_134, n_48, n_63, n_255, n_54, n_193, n_232, n_125, n_41, n_147, n_55, n_145, n_185, n_29, n_166, n_218, n_267, n_173, n_181, n_123, n_171, n_219, n_60, n_135, n_138, n_140, n_111, n_10, n_212, n_30, n_13, n_254, n_92, n_75, n_82, n_53, n_183, n_64, n_132, n_69, n_196, n_213, n_175, n_248, n_127, n_128, n_170, n_83, n_200, n_158, n_205, n_23, n_0, n_126, n_258, n_110, n_249, n_262, n_234, n_184, n_182, n_269, n_119, n_265, n_57, n_51, n_144, n_106, n_186, n_45, n_42, n_21, n_137, n_236, n_131, n_86, n_27, n_124, n_89, n_177, n_28, n_79, n_129, n_164, n_49, n_206, n_14, n_31, n_951, n_953);
input n_120;
input n_136;
input n_260;
input n_155;
input n_107;
input n_103;
input n_157;
input n_52;
input n_162;
input n_114;
input n_156;
input n_154;
input n_50;
input n_7;
input n_239;
input n_222;
input n_253;
input n_3;
input n_34;
input n_142;
input n_231;
input n_25;
input n_9;
input n_163;
input n_96;
input n_204;
input n_72;
input n_77;
input n_90;
input n_169;
input n_178;
input n_214;
input n_227;
input n_180;
input n_250;
input n_99;
input n_43;
input n_73;
input n_190;
input n_62;
input n_167;
input n_97;
input n_229;
input n_133;
input n_199;
input n_268;
input n_33;
input n_192;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_189;
input n_216;
input n_153;
input n_187;
input n_226;
input n_66;
input n_88;
input n_46;
input n_121;
input n_174;
input n_240;
input n_188;
input n_108;
input n_161;
input n_37;
input n_122;
input n_165;
input n_224;
input n_18;
input n_247;
input n_65;
input n_87;
input n_207;
input n_5;
input n_197;
input n_81;
input n_211;
input n_85;
input n_112;
input n_215;
input n_264;
input n_102;
input n_172;
input n_47;
input n_109;
input n_198;
input n_1;
input n_201;
input n_16;
input n_78;
input n_95;
input n_217;
input n_40;
input n_68;
input n_105;
input n_210;
input n_251;
input n_36;
input n_228;
input n_259;
input n_11;
input n_244;
input n_115;
input n_270;
input n_225;
input n_179;
input n_208;
input n_237;
input n_252;
input n_15;
input n_168;
input n_271;
input n_139;
input n_152;
input n_151;
input n_71;
input n_117;
input n_238;
input n_176;
input n_70;
input n_256;
input n_94;
input n_2;
input n_194;
input n_17;
input n_221;
input n_58;
input n_195;
input n_113;
input n_242;
input n_209;
input n_241;
input n_20;
input n_84;
input n_130;
input n_266;
input n_12;
input n_56;
input n_80;
input n_223;
input n_67;
input n_116;
input n_22;
input n_118;
input n_19;
input n_233;
input n_257;
input n_202;
input n_26;
input n_203;
input n_261;
input n_243;
input n_39;
input n_101;
input n_98;
input n_150;
input n_220;
input n_235;
input n_38;
input n_230;
input n_245;
input n_104;
input n_100;
input n_159;
input n_24;
input n_141;
input n_35;
input n_91;
input n_146;
input n_160;
input n_32;
input n_148;
input n_149;
input n_246;
input n_263;
input n_93;
input n_191;
input n_143;
input n_134;
input n_48;
input n_63;
input n_255;
input n_54;
input n_193;
input n_232;
input n_125;
input n_41;
input n_147;
input n_55;
input n_145;
input n_185;
input n_29;
input n_166;
input n_218;
input n_267;
input n_173;
input n_181;
input n_123;
input n_171;
input n_219;
input n_60;
input n_135;
input n_138;
input n_140;
input n_111;
input n_10;
input n_212;
input n_30;
input n_13;
input n_254;
input n_92;
input n_75;
input n_82;
input n_53;
input n_183;
input n_64;
input n_132;
input n_69;
input n_196;
input n_213;
input n_175;
input n_248;
input n_127;
input n_128;
input n_170;
input n_83;
input n_200;
input n_158;
input n_205;
input n_23;
input n_0;
input n_126;
input n_258;
input n_110;
input n_249;
input n_262;
input n_234;
input n_184;
input n_182;
input n_269;
input n_119;
input n_265;
input n_57;
input n_51;
input n_144;
input n_106;
input n_186;
input n_45;
input n_42;
input n_21;
input n_137;
input n_236;
input n_131;
input n_86;
input n_27;
input n_124;
input n_89;
input n_177;
input n_28;
input n_79;
input n_129;
input n_164;
input n_49;
input n_206;
input n_14;
input n_31;
output n_951;
output n_953;
wire n_890;
wire n_646;
wire n_107;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_239;
wire n_154;
wire n_7;
wire n_309;
wire n_944;
wire n_356;
wire n_895;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_929;
wire n_169;
wire n_370;
wire n_439;
wire n_384;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_44;
wire n_394;
wire n_189;
wire n_681;
wire n_226;
wire n_447;
wire n_352;
wire n_66;
wire n_379;
wire n_903;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_952;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_949;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_942;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_753;
wire n_176;
wire n_859;
wire n_438;
wire n_900;
wire n_869;
wire n_931;
wire n_935;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_838;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_410;
wire n_353;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_340;
wire n_301;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_555;
wire n_553;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_397;
wire n_315;
wire n_53;
wire n_880;
wire n_213;
wire n_797;
wire n_293;
wire n_836;
wire n_196;
wire n_312;
wire n_127;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_392;
wire n_120;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_816;
wire n_789;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_442;
wire n_324;
wire n_133;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_928;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_912;
wire n_920;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_905;
wire n_109;
wire n_332;
wire n_386;
wire n_934;
wire n_198;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_270;
wire n_115;
wire n_476;
wire n_765;
wire n_829;
wire n_599;
wire n_849;
wire n_715;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_911;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_800;
wire n_491;
wire n_711;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_906;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_879;
wire n_888;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_909;
wire n_493;
wire n_274;
wire n_910;
wire n_235;
wire n_150;
wire n_690;
wire n_533;
wire n_38;
wire n_272;
wire n_686;
wire n_100;
wire n_299;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_878;
wire n_812;
wire n_783;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_638;
wire n_171;
wire n_873;
wire n_899;
wire n_450;
wire n_585;
wire n_644;
wire n_140;
wire n_111;
wire n_779;
wire n_746;
wire n_212;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_704;
wire n_435;
wire n_728;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_921;
wire n_119;
wire n_667;
wire n_503;
wire n_856;
wire n_927;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_904;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_951;
wire n_348;
wire n_163;
wire n_96;
wire n_669;
wire n_685;
wire n_90;
wire n_72;
wire n_77;
wire n_594;
wire n_762;
wire n_214;
wire n_787;
wire n_740;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_908;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_946;
wire n_121;
wire n_286;
wire n_408;
wire n_206;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_537;
wire n_65;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_932;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_276;
wire n_297;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_815;
wire n_523;
wire n_854;
wire n_901;
wire n_528;
wire n_419;
wire n_252;
wire n_922;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_693;
wire n_785;
wire n_896;
wire n_739;
wire n_94;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_554;
wire n_597;
wire n_741;
wire n_705;
wire n_257;
wire n_698;
wire n_828;
wire n_722;
wire n_26;
wire n_203;
wire n_477;
wire n_460;
wire n_318;
wire n_243;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_337;
wire n_146;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_872;
wire n_539;
wire n_93;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_923;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_918;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_948;
wire n_732;
wire n_926;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_925;
wire n_915;
wire n_158;
wire n_205;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_89;
wire n_480;
wire n_939;
wire n_940;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_891;
wire n_580;
wire n_610;
wire n_938;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_34;
wire n_142;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_454;
wire n_395;
wire n_943;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_606;
wire n_190;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_565;
wire n_323;
wire n_59;
wire n_781;
wire n_914;
wire n_945;
wire n_852;
wire n_376;
wire n_902;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_88;
wire n_568;
wire n_46;
wire n_807;
wire n_717;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_87;
wire n_466;
wire n_207;
wire n_197;
wire n_541;
wire n_572;
wire n_81;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_919;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_416;
wire n_36;
wire n_916;
wire n_870;
wire n_889;
wire n_432;
wire n_913;
wire n_917;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_469;
wire n_369;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_520;
wire n_15;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_796;
wire n_804;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_907;
wire n_591;
wire n_391;
wire n_241;
wire n_209;
wire n_874;
wire n_20;
wire n_84;
wire n_782;
wire n_449;
wire n_832;
wire n_56;
wire n_412;
wire n_12;
wire n_455;
wire n_504;
wire n_67;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_930;
wire n_39;
wire n_101;
wire n_941;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_933;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_490;
wire n_472;
wire n_540;
wire n_947;
wire n_840;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_60;
wire n_138;
wire n_937;
wire n_936;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_924;
wire n_745;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_92;
wire n_313;
wire n_333;
wire n_358;
wire n_627;
wire n_706;
wire n_750;
wire n_589;
wire n_175;
wire n_897;
wire n_128;
wire n_415;
wire n_306;
wire n_31;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_625;
wire n_403;
wire n_144;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_436;
wire n_349;
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_199), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_252), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_56), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g275 ( .A(n_182), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_257), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_39), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_254), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_229), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_114), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_141), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_121), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_258), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_7), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_235), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_71), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_234), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_103), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_219), .Y(n_292) );
CKINVDCx16_ASAP7_75t_R g293 ( .A(n_216), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_245), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_161), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_94), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_118), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_109), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_261), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_255), .Y(n_300) );
INVx4_ASAP7_75t_R g301 ( .A(n_187), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_226), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_178), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_136), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_157), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_134), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_145), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_207), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_241), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_125), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_116), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_128), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_87), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_5), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_149), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_225), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_177), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_270), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_197), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_131), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_185), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_45), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_113), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_112), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_99), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_195), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_215), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_68), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_179), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_88), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_62), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_135), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_249), .B(n_256), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_92), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_239), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_183), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_231), .B(n_206), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_16), .B(n_243), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_189), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_180), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_269), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_236), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_137), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_248), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_30), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_194), .B(n_253), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_24), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_78), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_247), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_73), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_11), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_227), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_224), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_201), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_210), .Y(n_358) );
BUFx10_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_19), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_101), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_214), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_218), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_237), .Y(n_364) );
BUFx8_ASAP7_75t_SL g365 ( .A(n_147), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_100), .Y(n_366) );
BUFx2_ASAP7_75t_SL g367 ( .A(n_11), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_60), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_246), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_34), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_222), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_251), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_238), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_250), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_244), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_153), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_57), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_25), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_191), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_154), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_89), .Y(n_381) );
INVxp33_ASAP7_75t_SL g382 ( .A(n_223), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_90), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_33), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_51), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_44), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_167), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_150), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_64), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_232), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_61), .B(n_104), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_268), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_240), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_230), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_204), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_260), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_108), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_192), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_169), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_220), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_5), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_228), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_80), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_208), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_233), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_6), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_277), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_327), .B(n_0), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_399), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_293), .B(n_0), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_407), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_334), .B(n_1), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_334), .B(n_1), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_406), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_402), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_316), .Y(n_418) );
INVx5_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_406), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_374), .B(n_2), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_362), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_359), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_294), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_274), .A2(n_14), .B(n_13), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_310), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_430), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_413), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_408), .B(n_275), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_427), .B(n_336), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_415), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_410), .B(n_305), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g440 ( .A1(n_411), .A2(n_281), .B(n_278), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_414), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_416), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_426), .B(n_305), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_418), .B(n_414), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_412), .B(n_419), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_419), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_419), .B(n_354), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_428), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_432), .B(n_424), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_433), .B(n_425), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_434), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_441), .A2(n_423), .B1(n_409), .B2(n_382), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_440), .A2(n_417), .B1(n_367), .B2(n_397), .C(n_299), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_434), .B(n_272), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_448), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_439), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_446), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_442), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_444), .B(n_348), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_437), .B(n_273), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_435), .B(n_348), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_443), .B(n_284), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_445), .A2(n_292), .B1(n_314), .B2(n_276), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_447), .B(n_279), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_438), .B(n_282), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_436), .B(n_285), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_436), .B(n_286), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_449), .A2(n_361), .B1(n_378), .B2(n_343), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_453), .B(n_289), .C(n_287), .Y(n_472) );
OAI22x1_ASAP7_75t_L g473 ( .A1(n_463), .A2(n_336), .B1(n_365), .B2(n_429), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_466), .B(n_283), .Y(n_474) );
AOI21x1_ASAP7_75t_L g475 ( .A1(n_457), .A2(n_429), .B(n_391), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_450), .A2(n_291), .B(n_296), .C(n_295), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_460), .A2(n_303), .B(n_298), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_451), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_455), .Y(n_479) );
NOR2x1p5_ASAP7_75t_SL g480 ( .A(n_464), .B(n_340), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_469), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_460), .B(n_288), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_452), .B(n_290), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_454), .A2(n_308), .B(n_306), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_462), .B(n_297), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_461), .A2(n_462), .B(n_459), .Y(n_488) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_461), .B(n_312), .C(n_311), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_455), .A2(n_349), .B1(n_315), .B2(n_317), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_468), .A2(n_318), .B(n_313), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_468), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_465), .A2(n_467), .B(n_470), .Y(n_493) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_468), .A2(n_422), .A3(n_420), .B1(n_415), .B2(n_364), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_482), .Y(n_495) );
OAI21x1_ASAP7_75t_L g496 ( .A1(n_475), .A2(n_321), .B(n_320), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_479), .Y(n_497) );
OAI21x1_ASAP7_75t_L g498 ( .A1(n_493), .A2(n_325), .B(n_322), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_485), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_300), .B1(n_304), .B2(n_302), .Y(n_500) );
AOI21xp5_ASAP7_75t_SL g501 ( .A1(n_473), .A2(n_307), .B(n_280), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_471), .B(n_309), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_488), .A2(n_331), .B(n_326), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_479), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_491), .A2(n_333), .B(n_332), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_486), .A2(n_337), .B(n_335), .Y(n_508) );
AOI21x1_ASAP7_75t_SL g509 ( .A1(n_487), .A2(n_301), .B(n_328), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_479), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_477), .A2(n_350), .B(n_345), .Y(n_511) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_490), .A2(n_363), .B(n_356), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_472), .B(n_7), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_484), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_483), .A2(n_323), .B1(n_324), .B2(n_319), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_476), .B(n_329), .Y(n_516) );
AOI21x1_ASAP7_75t_L g517 ( .A1(n_474), .A2(n_376), .B(n_373), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_489), .B(n_330), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_480), .B(n_339), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_494), .Y(n_520) );
BUFx4_ASAP7_75t_SL g521 ( .A(n_494), .Y(n_521) );
CKINVDCx8_ASAP7_75t_R g522 ( .A(n_494), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_488), .A2(n_380), .B(n_377), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_488), .A2(n_385), .B(n_383), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_499), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_506), .B(n_8), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_502), .Y(n_528) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_496), .A2(n_372), .B(n_338), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_514), .B(n_8), .Y(n_530) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_520), .A2(n_398), .B(n_386), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_503), .A2(n_401), .B1(n_403), .B2(n_400), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_513), .B(n_9), .Y(n_533) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_498), .A2(n_387), .B(n_381), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_505), .B(n_9), .Y(n_535) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_509), .A2(n_405), .B(n_388), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_512), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_507), .A2(n_404), .B1(n_389), .B2(n_346), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_517), .Y(n_539) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_524), .A2(n_341), .B(n_17), .Y(n_540) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_504), .A2(n_18), .B(n_15), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_505), .B(n_10), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_523), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_508), .A2(n_422), .B(n_420), .Y(n_544) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_507), .A2(n_344), .B(n_342), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_510), .A2(n_21), .B(n_20), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_516), .B(n_10), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_497), .Y(n_549) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_511), .A2(n_351), .B(n_347), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_503), .B(n_12), .Y(n_552) );
AOI22x1_ASAP7_75t_L g553 ( .A1(n_501), .A2(n_395), .B1(n_394), .B2(n_393), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_519), .A2(n_353), .B(n_352), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_518), .A2(n_357), .B(n_355), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_521), .B(n_12), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_522), .B(n_22), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_515), .A2(n_360), .B(n_358), .Y(n_559) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_520), .A2(n_23), .B(n_26), .Y(n_560) );
CKINVDCx14_ASAP7_75t_R g561 ( .A(n_499), .Y(n_561) );
NOR2xp33_ASAP7_75t_SL g562 ( .A(n_503), .B(n_366), .Y(n_562) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_520), .A2(n_27), .B(n_28), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_499), .B(n_368), .Y(n_564) );
AOI21xp33_ASAP7_75t_L g565 ( .A1(n_519), .A2(n_370), .B(n_369), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_514), .B(n_371), .Y(n_566) );
OAI21x1_ASAP7_75t_L g567 ( .A1(n_496), .A2(n_29), .B(n_31), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_503), .A2(n_392), .B1(n_390), .B2(n_384), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_524), .A2(n_375), .B(n_35), .C(n_36), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_495), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_528), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_546), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_525), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_546), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_561), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_531), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_570), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_571), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_543), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_551), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_527), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_539), .B(n_32), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_535), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_549), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_549), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_530), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_37), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_548), .A2(n_38), .B(n_40), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_567), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_552), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_556), .B(n_566), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_558), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_538), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_550), .Y(n_600) );
OA21x2_ASAP7_75t_L g601 ( .A1(n_534), .A2(n_529), .B(n_540), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_569), .A2(n_41), .B(n_42), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
AO21x1_ASAP7_75t_SL g604 ( .A1(n_532), .A2(n_43), .B(n_46), .Y(n_604) );
NOR2xp33_ASAP7_75t_SL g605 ( .A(n_557), .B(n_47), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_550), .Y(n_606) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_544), .A2(n_563), .B(n_560), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_545), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
AOI21x1_ASAP7_75t_L g610 ( .A1(n_557), .A2(n_48), .B(n_49), .Y(n_610) );
AO21x2_ASAP7_75t_L g611 ( .A1(n_541), .A2(n_50), .B(n_52), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_555), .Y(n_614) );
BUFx2_ASAP7_75t_SL g615 ( .A(n_553), .Y(n_615) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_554), .A2(n_53), .B(n_54), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_559), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_568), .B(n_55), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
INVx3_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
OAI21x1_ASAP7_75t_L g623 ( .A1(n_529), .A2(n_58), .B(n_59), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_537), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_526), .B(n_271), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_526), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_546), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_526), .B(n_63), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_528), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_528), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_526), .B(n_65), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_528), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_528), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_526), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_528), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_546), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_528), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_526), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_526), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_528), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_526), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_526), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_528), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_546), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_526), .B(n_66), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_537), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_528), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_526), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_626), .B(n_67), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_583), .B(n_69), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_605), .A2(n_70), .B1(n_72), .B2(n_74), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_582), .B(n_75), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_634), .B(n_76), .Y(n_656) );
INVx2_ASAP7_75t_SL g657 ( .A(n_578), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_629), .Y(n_658) );
OA21x2_ASAP7_75t_L g659 ( .A1(n_595), .A2(n_77), .B(n_79), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_582), .B(n_81), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_638), .B(n_82), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_574), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_630), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_632), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_598), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_633), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_635), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_637), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_575), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_639), .B(n_83), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_640), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_642), .B(n_84), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_649), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_575), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_605), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_612), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_585), .B(n_85), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_643), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_648), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_576), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_588), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_577), .Y(n_683) );
INVx4_ASAP7_75t_L g684 ( .A(n_644), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_585), .B(n_86), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_620), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_597), .B(n_91), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_583), .B(n_93), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_650), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_581), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_599), .B(n_95), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_587), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_591), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_589), .B(n_267), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_592), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_619), .B(n_96), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_576), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_596), .B(n_265), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_613), .B(n_97), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_573), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_624), .B(n_98), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_584), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_584), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_573), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_624), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_646), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_617), .B(n_102), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_622), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_646), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_631), .B(n_645), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_614), .B(n_105), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_593), .B(n_106), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_622), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_625), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_628), .B(n_107), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_627), .B(n_110), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_627), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_620), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_610), .A2(n_111), .B1(n_115), .B2(n_117), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_636), .B(n_119), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_647), .B(n_263), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_644), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_644), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_636), .B(n_120), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_621), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_621), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_647), .B(n_122), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_579), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_600), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_608), .B(n_123), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_579), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_580), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_609), .B(n_124), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_580), .B(n_126), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_606), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_586), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_586), .Y(n_737) );
BUFx2_ASAP7_75t_L g738 ( .A(n_594), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_616), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_618), .B(n_127), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_623), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_611), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_604), .B(n_129), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_594), .B(n_130), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_590), .B(n_132), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_672), .B(n_607), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_735), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_695), .B(n_607), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_683), .B(n_602), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_674), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_657), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_682), .B(n_601), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_726), .B(n_603), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_690), .B(n_602), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_654), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_692), .B(n_601), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_658), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_669), .Y(n_758) );
NOR2x1p5_ASAP7_75t_L g759 ( .A(n_681), .B(n_615), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_693), .B(n_611), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_663), .B(n_133), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_664), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_669), .B(n_138), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_666), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_667), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_675), .B(n_139), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_686), .B(n_140), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_668), .B(n_142), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_671), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_679), .B(n_143), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_705), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_706), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_680), .B(n_144), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_689), .B(n_146), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_665), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_686), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_665), .Y(n_778) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_722), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_714), .B(n_704), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_718), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_725), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_702), .B(n_148), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_736), .B(n_151), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_709), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_708), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_703), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_713), .B(n_152), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_717), .B(n_155), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_737), .B(n_156), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_729), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_710), .B(n_158), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_728), .Y(n_793) );
INVx1_ASAP7_75t_SL g794 ( .A(n_677), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_731), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_732), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_701), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_681), .B(n_159), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_723), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_684), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_697), .B(n_160), .Y(n_801) );
CKINVDCx16_ASAP7_75t_R g802 ( .A(n_662), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_684), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_697), .B(n_162), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_687), .B(n_163), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_678), .B(n_164), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_741), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_700), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_685), .B(n_165), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_676), .B(n_166), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_696), .B(n_168), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_701), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_676), .B(n_170), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_699), .B(n_171), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_738), .B(n_172), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_780), .B(n_739), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_781), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_758), .B(n_655), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_776), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_799), .B(n_739), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_765), .B(n_660), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_802), .B(n_712), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_795), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_786), .B(n_743), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_791), .B(n_742), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_757), .B(n_651), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_778), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_762), .B(n_656), .Y(n_828) );
AND2x4_ASAP7_75t_SL g829 ( .A(n_808), .B(n_716), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_759), .B(n_720), .Y(n_830) );
INVx1_ASAP7_75t_SL g831 ( .A(n_779), .Y(n_831) );
NOR2x1p5_ASAP7_75t_L g832 ( .A(n_800), .B(n_698), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_750), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_764), .B(n_661), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_777), .B(n_734), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_755), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_766), .B(n_670), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_746), .B(n_724), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_770), .B(n_673), .Y(n_839) );
BUFx2_ASAP7_75t_L g840 ( .A(n_779), .Y(n_840) );
INVxp67_ASAP7_75t_L g841 ( .A(n_748), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_747), .B(n_691), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_803), .B(n_653), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_747), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_796), .B(n_691), .Y(n_845) );
INVxp33_ASAP7_75t_L g846 ( .A(n_779), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_782), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_793), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_751), .B(n_711), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_793), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_772), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_785), .Y(n_852) );
NAND2xp33_ASAP7_75t_L g853 ( .A(n_794), .B(n_744), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_772), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_773), .Y(n_855) );
NOR2xp33_ASAP7_75t_R g856 ( .A(n_805), .B(n_727), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_773), .Y(n_857) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_752), .Y(n_858) );
OR2x6_ASAP7_75t_L g859 ( .A(n_830), .B(n_763), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_853), .A2(n_792), .B1(n_797), .B2(n_812), .Y(n_860) );
OR2x6_ASAP7_75t_L g861 ( .A(n_830), .B(n_763), .Y(n_861) );
INVx3_ASAP7_75t_L g862 ( .A(n_829), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_836), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_817), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_843), .B(n_760), .C(n_815), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_844), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_858), .Y(n_867) );
AND2x4_ASAP7_75t_L g868 ( .A(n_820), .B(n_756), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_816), .B(n_807), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_824), .B(n_753), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_822), .B(n_810), .Y(n_871) );
INVxp67_ASAP7_75t_L g872 ( .A(n_840), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_838), .B(n_753), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_819), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_827), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_838), .B(n_787), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_841), .B(n_807), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_847), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_851), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_833), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_848), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_850), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_841), .B(n_812), .Y(n_883) );
INVx2_ASAP7_75t_SL g884 ( .A(n_831), .Y(n_884) );
INVxp67_ASAP7_75t_L g885 ( .A(n_849), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_867), .B(n_825), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_865), .B(n_843), .C(n_852), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_864), .Y(n_888) );
OAI322xp33_ASAP7_75t_L g889 ( .A1(n_883), .A2(n_821), .A3(n_818), .B1(n_835), .B2(n_845), .C1(n_842), .C2(n_854), .Y(n_889) );
NAND2x2_ASAP7_75t_L g890 ( .A(n_884), .B(n_832), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_880), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_879), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_859), .A2(n_846), .B1(n_831), .B2(n_813), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_859), .A2(n_839), .B1(n_828), .B2(n_826), .Y(n_894) );
AOI322xp5_ASAP7_75t_L g895 ( .A1(n_871), .A2(n_834), .A3(n_837), .B1(n_842), .B2(n_845), .C1(n_857), .C2(n_855), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_861), .A2(n_767), .B1(n_768), .B2(n_823), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_877), .B(n_749), .Y(n_897) );
NAND2xp33_ASAP7_75t_SL g898 ( .A(n_862), .B(n_856), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g899 ( .A(n_860), .B(n_767), .Y(n_899) );
NAND2x1p5_ASAP7_75t_L g900 ( .A(n_873), .B(n_768), .Y(n_900) );
INVx1_ASAP7_75t_SL g901 ( .A(n_870), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_868), .B(n_754), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_895), .B(n_874), .Y(n_903) );
INVxp67_ASAP7_75t_L g904 ( .A(n_898), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_890), .A2(n_861), .B1(n_876), .B2(n_869), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_887), .B(n_872), .C(n_875), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_888), .Y(n_907) );
OAI21xp33_ASAP7_75t_SL g908 ( .A1(n_899), .A2(n_885), .B(n_878), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_897), .B(n_863), .C(n_881), .Y(n_909) );
AOI222xp33_ASAP7_75t_L g910 ( .A1(n_886), .A2(n_882), .B1(n_866), .B2(n_869), .C1(n_868), .C2(n_775), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_892), .Y(n_911) );
AOI32xp33_ASAP7_75t_L g912 ( .A1(n_893), .A2(n_809), .A3(n_788), .B1(n_789), .B2(n_814), .Y(n_912) );
O2A1O1Ixp5_ASAP7_75t_L g913 ( .A1(n_889), .A2(n_798), .B(n_804), .C(n_784), .Y(n_913) );
OAI21xp5_ASAP7_75t_SL g914 ( .A1(n_896), .A2(n_811), .B(n_740), .Y(n_914) );
OAI21xp33_ASAP7_75t_L g915 ( .A1(n_908), .A2(n_894), .B(n_902), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_904), .A2(n_901), .B(n_894), .Y(n_916) );
AOI211xp5_ASAP7_75t_SL g917 ( .A1(n_903), .A2(n_719), .B(n_801), .C(n_721), .Y(n_917) );
OAI21xp33_ASAP7_75t_L g918 ( .A1(n_910), .A2(n_900), .B(n_891), .Y(n_918) );
AOI211xp5_ASAP7_75t_L g919 ( .A1(n_914), .A2(n_719), .B(n_769), .C(n_806), .Y(n_919) );
AOI221x1_ASAP7_75t_L g920 ( .A1(n_906), .A2(n_774), .B1(n_790), .B2(n_783), .C(n_771), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_905), .B(n_761), .Y(n_921) );
NOR2xp67_ASAP7_75t_L g922 ( .A(n_909), .B(n_173), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_915), .A2(n_913), .B1(n_912), .B2(n_907), .C(n_911), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_916), .Y(n_924) );
NOR2x1_ASAP7_75t_L g925 ( .A(n_922), .B(n_715), .Y(n_925) );
NOR3xp33_ASAP7_75t_L g926 ( .A(n_918), .B(n_652), .C(n_688), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_921), .B(n_694), .Y(n_927) );
NOR3xp33_ASAP7_75t_L g928 ( .A(n_924), .B(n_919), .C(n_917), .Y(n_928) );
NAND4xp25_ASAP7_75t_SL g929 ( .A(n_923), .B(n_920), .C(n_652), .D(n_688), .Y(n_929) );
NAND3x2_ASAP7_75t_L g930 ( .A(n_926), .B(n_707), .C(n_176), .Y(n_930) );
NAND4xp25_ASAP7_75t_SL g931 ( .A(n_925), .B(n_733), .C(n_730), .D(n_745), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_929), .B(n_927), .Y(n_932) );
CKINVDCx16_ASAP7_75t_R g933 ( .A(n_928), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_930), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_931), .B(n_659), .Y(n_935) );
NAND2x1p5_ASAP7_75t_L g936 ( .A(n_934), .B(n_659), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_933), .Y(n_937) );
BUFx3_ASAP7_75t_L g938 ( .A(n_932), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_937), .A2(n_935), .B1(n_733), .B2(n_730), .Y(n_939) );
NAND2x1p5_ASAP7_75t_L g940 ( .A(n_938), .B(n_745), .Y(n_940) );
OR2x6_ASAP7_75t_L g941 ( .A(n_936), .B(n_174), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_939), .B(n_181), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_940), .B(n_184), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_941), .B(n_186), .Y(n_944) );
AO21x2_ASAP7_75t_L g945 ( .A1(n_942), .A2(n_188), .B(n_190), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_943), .B(n_193), .Y(n_946) );
OAI21xp5_ASAP7_75t_L g947 ( .A1(n_946), .A2(n_944), .B(n_198), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_945), .A2(n_196), .B(n_200), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_948), .B(n_202), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_947), .A2(n_203), .B1(n_205), .B2(n_209), .Y(n_950) );
UNKNOWN g951 ( );
OR2x6_ASAP7_75t_L g952 ( .A(n_949), .B(n_211), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_951), .A2(n_952), .B1(n_212), .B2(n_213), .Y(n_953) );
endmodule