module fake_ariane_1831_n_1174 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1174);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1174;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_908;
wire n_850;
wire n_788;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_905;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_1134;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_1099;
wire n_928;
wire n_271;
wire n_1153;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_1080;
wire n_899;
wire n_1148;
wire n_576;
wire n_843;
wire n_920;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_543;
wire n_362;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_772;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_1110;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_118),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_6),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_134),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_18),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_52),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_170),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_79),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_67),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_65),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_177),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_92),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_83),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_47),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_129),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_75),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_46),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_85),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_96),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_25),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_148),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_208),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_132),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_93),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_213),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_95),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_159),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_68),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_113),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_137),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_128),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_73),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_62),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_10),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_71),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_237),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_280),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_255),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_223),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_276),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_0),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_271),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_241),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_241),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_241),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_223),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_229),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_258),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_279),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_256),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_322),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_260),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_260),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_258),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_220),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_221),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_225),
.Y(n_355)
);

OAI21x1_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_230),
.B(n_226),
.Y(n_356)
);

CKINVDCx11_ASAP7_75t_R g357 ( 
.A(n_336),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_231),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_305),
.A2(n_272),
.B1(n_282),
.B2(n_287),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_302),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_319),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_272),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_299),
.A2(n_235),
.B(n_233),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_242),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_321),
.B(n_282),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_287),
.B1(n_289),
.B2(n_288),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_334),
.A2(n_291),
.B1(n_286),
.B2(n_285),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

AND2x2_ASAP7_75t_SL g387 ( 
.A(n_324),
.B(n_38),
.Y(n_387)
);

CKINVDCx11_ASAP7_75t_R g388 ( 
.A(n_336),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_326),
.B(n_246),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_247),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_248),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_343),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_382),
.B(n_303),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_361),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_382),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_372),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_372),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_342),
.B(n_293),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_355),
.B(n_293),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_372),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_361),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_378),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_378),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_347),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_383),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_383),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_342),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_376),
.B(n_316),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_377),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_359),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_375),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_391),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_381),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_351),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_346),
.B(n_311),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_354),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_348),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_348),
.B(n_314),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_348),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_368),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_389),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_348),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_344),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_344),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_344),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_344),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_344),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_368),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_376),
.B(n_316),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_392),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_376),
.B(n_295),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_392),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_365),
.B(n_310),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_344),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_344),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_368),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_365),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_387),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_443),
.B(n_387),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_445),
.B(n_387),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_341),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_429),
.B(n_330),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_397),
.B(n_386),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_368),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_386),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_386),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_294),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_433),
.B(n_390),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_390),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_390),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_413),
.B(n_380),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_296),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_390),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_368),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_368),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_368),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_403),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_464),
.B(n_379),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_463),
.B(n_376),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_415),
.B(n_379),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_469),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_401),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_379),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_423),
.A2(n_424),
.B1(n_418),
.B2(n_420),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_434),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g523 ( 
.A(n_423),
.B(n_340),
.C(n_332),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_385),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_439),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_469),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_419),
.B(n_385),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_460),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_459),
.A2(n_298),
.B1(n_308),
.B2(n_292),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_456),
.B(n_308),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_407),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_417),
.B(n_296),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_444),
.B(n_394),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_369),
.C(n_385),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_466),
.B(n_393),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_452),
.B(n_393),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_410),
.B(n_309),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_466),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_428),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_474),
.B(n_453),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_428),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

NOR3xp33_ASAP7_75t_L g561 ( 
.A(n_477),
.B(n_414),
.C(n_412),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_416),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_511),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_506),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_498),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_475),
.A2(n_420),
.B1(n_406),
.B2(n_455),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_474),
.B(n_465),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_513),
.B(n_406),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_476),
.A2(n_307),
.B1(n_304),
.B2(n_370),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_538),
.B(n_370),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_489),
.B(n_393),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_493),
.B(n_489),
.C(n_478),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_395),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_481),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_466),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_373),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_487),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_497),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_551),
.B(n_356),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_521),
.A2(n_307),
.B1(n_257),
.B2(n_259),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_532),
.B(n_373),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_551),
.B(n_356),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_523),
.A2(n_350),
.B1(n_353),
.B2(n_369),
.C(n_371),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_395),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_508),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_541),
.B(n_350),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_492),
.B(n_353),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_520),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_522),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_512),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_530),
.B(n_369),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_480),
.B(n_369),
.C(n_395),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_515),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_534),
.B(n_371),
.C(n_263),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_492),
.B(n_371),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_556),
.B(n_264),
.C(n_254),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_501),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_509),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_552),
.B(n_371),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_394),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_536),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_479),
.B(n_394),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_505),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_530),
.B(n_394),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_479),
.B(n_371),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_492),
.B(n_371),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_556),
.B(n_269),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_507),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_507),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_518),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_526),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_333),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_598),
.A2(n_542),
.B(n_484),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_598),
.A2(n_472),
.B1(n_471),
.B2(n_482),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_492),
.Y(n_629)
);

NOR2x1p5_ASAP7_75t_SL g630 ( 
.A(n_622),
.B(n_623),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_557),
.B(n_510),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_600),
.B(n_555),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_609),
.B(n_498),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_612),
.A2(n_524),
.B(n_484),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_L g636 ( 
.A1(n_619),
.A2(n_537),
.B(n_539),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_612),
.A2(n_550),
.B(n_502),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_523),
.B(n_504),
.C(n_505),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_585),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_582),
.A2(n_580),
.B(n_578),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_564),
.B(n_510),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_570),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_578),
.A2(n_550),
.B(n_502),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_559),
.B(n_548),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_L g645 ( 
.A1(n_616),
.A2(n_553),
.B(n_549),
.Y(n_645)
);

BUFx4f_ASAP7_75t_L g646 ( 
.A(n_566),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_SL g647 ( 
.A1(n_586),
.A2(n_472),
.B(n_504),
.C(n_518),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_571),
.A2(n_503),
.B1(n_535),
.B2(n_541),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_568),
.B(n_510),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_603),
.A2(n_503),
.B(n_535),
.C(n_545),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_575),
.B(n_510),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_575),
.B(n_534),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_611),
.B(n_494),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_604),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_561),
.B(n_543),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_614),
.A2(n_545),
.B(n_529),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_572),
.B(n_494),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_610),
.B(n_613),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_494),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_580),
.A2(n_554),
.B(n_516),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_608),
.B(n_529),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_614),
.A2(n_531),
.B(n_500),
.Y(n_663)
);

NOR3xp33_ASAP7_75t_L g664 ( 
.A(n_606),
.B(n_500),
.C(n_275),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_608),
.A2(n_531),
.B1(n_544),
.B2(n_546),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_592),
.A2(n_554),
.B(n_516),
.Y(n_666)
);

BUFx4f_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

CKINVDCx10_ASAP7_75t_R g668 ( 
.A(n_565),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_544),
.B1(n_546),
.B2(n_531),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_599),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_SL g672 ( 
.A1(n_558),
.A2(n_544),
.B(n_618),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_595),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_R g674 ( 
.A(n_624),
.B(n_495),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_617),
.A2(n_531),
.B(n_547),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_L g676 ( 
.A1(n_624),
.A2(n_277),
.B(n_274),
.Y(n_676)
);

OAI321xp33_ASAP7_75t_L g677 ( 
.A1(n_590),
.A2(n_517),
.A3(n_516),
.B1(n_495),
.B2(n_364),
.C(n_366),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_621),
.B(n_560),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_576),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_L g680 ( 
.A(n_588),
.B(n_546),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_626),
.A2(n_517),
.B(n_495),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_577),
.B(n_517),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_596),
.B(n_547),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_621),
.B(n_278),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_626),
.A2(n_547),
.B(n_284),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_597),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_558),
.A2(n_366),
.B(n_364),
.C(n_363),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_617),
.A2(n_547),
.B(n_362),
.Y(n_688)
);

CKINVDCx14_ASAP7_75t_R g689 ( 
.A(n_595),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_569),
.A2(n_362),
.B(n_345),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_583),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_589),
.A2(n_362),
.B(n_345),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_573),
.B(n_3),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_667),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_634),
.A2(n_601),
.B(n_590),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_674),
.Y(n_696)
);

NOR2x1_ASAP7_75t_SL g697 ( 
.A(n_651),
.B(n_563),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_659),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_667),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_637),
.A2(n_640),
.B(n_643),
.Y(n_700)
);

BUFx5_ASAP7_75t_L g701 ( 
.A(n_679),
.Y(n_701)
);

AOI33xp33_ASAP7_75t_L g702 ( 
.A1(n_644),
.A2(n_662),
.A3(n_686),
.B1(n_669),
.B2(n_636),
.B3(n_670),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_652),
.B(n_581),
.Y(n_703)
);

OR2x2_ASAP7_75t_SL g704 ( 
.A(n_658),
.B(n_615),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_645),
.A2(n_615),
.B1(n_584),
.B2(n_591),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_627),
.A2(n_573),
.B(n_615),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_668),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_660),
.A2(n_573),
.B1(n_567),
.B2(n_574),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_677),
.A2(n_594),
.B(n_593),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_654),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_642),
.B(n_625),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_649),
.A2(n_605),
.B1(n_602),
.B2(n_594),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_682),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_655),
.A2(n_632),
.B(n_693),
.C(n_638),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_654),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_SL g717 ( 
.A(n_633),
.B(n_4),
.C(n_5),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_677),
.A2(n_363),
.B(n_345),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_689),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_639),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_653),
.B(n_4),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_678),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_673),
.B(n_5),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_364),
.B1(n_363),
.B2(n_366),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_676),
.B(n_6),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_630),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_673),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_646),
.Y(n_728)
);

AO22x1_ASAP7_75t_L g729 ( 
.A1(n_664),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_646),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_648),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_671),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_629),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_733)
);

AOI21xp33_ASAP7_75t_L g734 ( 
.A1(n_631),
.A2(n_14),
.B(n_15),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_663),
.A2(n_40),
.B(n_39),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_654),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_657),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_657),
.B(n_15),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_657),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_641),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_675),
.A2(n_44),
.B(n_42),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_635),
.B(n_16),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_680),
.B(n_16),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_628),
.A2(n_17),
.B(n_18),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

CKINVDCx8_ASAP7_75t_R g746 ( 
.A(n_684),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_647),
.A2(n_17),
.B(n_19),
.C(n_20),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_672),
.B(n_20),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_691),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_691),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_665),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_650),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_683),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_753)
);

BUFx12f_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_681),
.B(n_45),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_692),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_656),
.B(n_26),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_698),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_736),
.Y(n_759)
);

BUFx2_ASAP7_75t_SL g760 ( 
.A(n_728),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_736),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_699),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_727),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_703),
.B(n_661),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_732),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_750),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_720),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_736),
.B(n_688),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_716),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_748),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_708),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_716),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_737),
.B(n_666),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_699),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_749),
.A2(n_685),
.B1(n_690),
.B2(n_29),
.Y(n_775)
);

INVx5_ASAP7_75t_SL g776 ( 
.A(n_748),
.Y(n_776)
);

BUFx2_ASAP7_75t_R g777 ( 
.A(n_739),
.Y(n_777)
);

BUFx12f_ASAP7_75t_L g778 ( 
.A(n_696),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_705),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_716),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_719),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_714),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_694),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_737),
.B(n_49),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_704),
.B(n_722),
.Y(n_785)
);

INVx5_ASAP7_75t_L g786 ( 
.A(n_694),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_737),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_730),
.B(n_27),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_711),
.Y(n_789)
);

INVx6_ASAP7_75t_SL g790 ( 
.A(n_746),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_711),
.B(n_50),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_712),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_738),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_751),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_751),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_701),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_745),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_743),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_754),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_701),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_756),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_701),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_756),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_717),
.Y(n_805)
);

BUFx5_ASAP7_75t_L g806 ( 
.A(n_740),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_701),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_28),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_757),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_707),
.B(n_709),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_756),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_715),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_697),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_742),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_726),
.B(n_28),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_706),
.B(n_29),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_702),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_744),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_755),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_733),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_752),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_713),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_741),
.B(n_51),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_695),
.B(n_30),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_747),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_731),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_710),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_700),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_753),
.B(n_31),
.Y(n_833)
);

INVx6_ASAP7_75t_L g834 ( 
.A(n_778),
.Y(n_834)
);

AO21x2_ASAP7_75t_L g835 ( 
.A1(n_810),
.A2(n_735),
.B(n_718),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_SL g836 ( 
.A1(n_819),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_828),
.A2(n_764),
.B(n_773),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_763),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_828),
.A2(n_724),
.B(n_140),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_764),
.A2(n_139),
.B(n_218),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_763),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_773),
.A2(n_138),
.B(n_217),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_813),
.B(n_35),
.C(n_36),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_814),
.A2(n_135),
.B(n_216),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_779),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_814),
.A2(n_133),
.B(n_215),
.Y(n_846)
);

CKINVDCx14_ASAP7_75t_R g847 ( 
.A(n_771),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_758),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_827),
.A2(n_131),
.B(n_212),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_782),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_829),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_770),
.B(n_53),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_832),
.A2(n_141),
.B(n_54),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_765),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_810),
.A2(n_37),
.B(n_219),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_803),
.A2(n_55),
.B(n_56),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_803),
.A2(n_57),
.B(n_59),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_797),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_795),
.A2(n_60),
.B(n_61),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_795),
.B(n_211),
.Y(n_860)
);

AOI222xp33_ASAP7_75t_L g861 ( 
.A1(n_823),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.C1(n_70),
.C2(n_72),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_807),
.A2(n_74),
.B(n_76),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_794),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_815),
.B(n_793),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_766),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_813),
.B(n_77),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_793),
.B(n_78),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_820),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_868)
);

AO31x2_ASAP7_75t_L g869 ( 
.A1(n_826),
.A2(n_84),
.A3(n_86),
.B(n_87),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_820),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_820),
.A2(n_94),
.B(n_97),
.C(n_99),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_781),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_792),
.B(n_100),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_794),
.B(n_101),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_799),
.A2(n_102),
.B(n_103),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_766),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_SL g877 ( 
.A1(n_833),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_877)
);

AO31x2_ASAP7_75t_L g878 ( 
.A1(n_801),
.A2(n_107),
.A3(n_108),
.B(n_109),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_796),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_809),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_802),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_812),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_830),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_883)
);

AO21x2_ASAP7_75t_L g884 ( 
.A1(n_824),
.A2(n_115),
.B(n_116),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_785),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_800),
.B(n_117),
.Y(n_886)
);

OAI221xp5_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.C(n_122),
.Y(n_887)
);

CKINVDCx6p67_ASAP7_75t_R g888 ( 
.A(n_760),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_SL g889 ( 
.A1(n_770),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_817),
.A2(n_130),
.B(n_142),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_833),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_891)
);

OAI21x1_ASAP7_75t_SL g892 ( 
.A1(n_821),
.A2(n_147),
.B(n_150),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_806),
.B(n_812),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_759),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_816),
.A2(n_151),
.B(n_152),
.C(n_153),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_791),
.A2(n_154),
.B(n_155),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_805),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_880),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_893),
.B(n_796),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_838),
.B(n_806),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_845),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_879),
.B(n_806),
.Y(n_902)
);

AO21x2_ASAP7_75t_L g903 ( 
.A1(n_835),
.A2(n_817),
.B(n_818),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_837),
.A2(n_840),
.B(n_839),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_880),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_854),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_850),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_848),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_865),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_876),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_894),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_885),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_882),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_879),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_838),
.B(n_825),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_861),
.A2(n_816),
.B1(n_798),
.B2(n_770),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_SL g917 ( 
.A1(n_866),
.A2(n_800),
.B(n_767),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_860),
.A2(n_768),
.B(n_808),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_841),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_853),
.A2(n_784),
.B(n_783),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_841),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_863),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_855),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_855),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_859),
.A2(n_783),
.B(n_774),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_858),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_835),
.A2(n_775),
.B(n_768),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_863),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_864),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_861),
.A2(n_776),
.B1(n_806),
.B2(n_831),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_894),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_860),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_887),
.A2(n_831),
.B1(n_786),
.B2(n_774),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_897),
.A2(n_776),
.B1(n_806),
.B2(n_831),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_874),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_878),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_866),
.B(n_804),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_834),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_881),
.Y(n_939)
);

BUFx2_ASAP7_75t_R g940 ( 
.A(n_872),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_873),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_867),
.B(n_878),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_890),
.A2(n_811),
.B(n_777),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_878),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_851),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_894),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_869),
.Y(n_947)
);

AO21x1_ASAP7_75t_SL g948 ( 
.A1(n_874),
.A2(n_811),
.B(n_777),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_R g949 ( 
.A(n_942),
.B(n_852),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_945),
.A2(n_897),
.B1(n_843),
.B2(n_887),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_915),
.B(n_888),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_907),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_929),
.B(n_834),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_898),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_905),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_919),
.B(n_834),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_921),
.B(n_886),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_942),
.A2(n_883),
.B1(n_891),
.B2(n_852),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_906),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_922),
.Y(n_960)
);

CKINVDCx16_ASAP7_75t_R g961 ( 
.A(n_901),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_922),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_906),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_915),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_908),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_907),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_912),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_901),
.B(n_847),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_902),
.B(n_852),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_938),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_940),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_922),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_909),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_939),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_914),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_926),
.Y(n_976)
);

AO21x2_ASAP7_75t_L g977 ( 
.A1(n_923),
.A2(n_892),
.B(n_871),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_SL g978 ( 
.A(n_917),
.B(n_788),
.C(n_851),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_910),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_914),
.B(n_769),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_933),
.A2(n_871),
.B(n_877),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_930),
.A2(n_891),
.B1(n_883),
.B2(n_889),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_938),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_L g984 ( 
.A(n_932),
.B(n_895),
.C(n_836),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_900),
.B(n_886),
.C(n_868),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_913),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_952),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_952),
.Y(n_988)
);

AOI221xp5_ASAP7_75t_L g989 ( 
.A1(n_950),
.A2(n_836),
.B1(n_923),
.B2(n_916),
.C(n_903),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_966),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_959),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_963),
.Y(n_992)
);

AND2x4_ASAP7_75t_SL g993 ( 
.A(n_969),
.B(n_937),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_954),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_955),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_966),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_960),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_973),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_964),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_979),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_981),
.A2(n_943),
.B(n_918),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_964),
.B(n_975),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_975),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_965),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_967),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_976),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_957),
.B(n_903),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_968),
.B(n_935),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_971),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_971),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_1009),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_993),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_991),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_993),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_1007),
.A2(n_978),
.B(n_950),
.C(n_958),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1008),
.B(n_953),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_991),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_992),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_987),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1006),
.B(n_957),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_999),
.B(n_970),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_1002),
.B(n_980),
.Y(n_1022)
);

AOI222xp33_ASAP7_75t_L g1023 ( 
.A1(n_989),
.A2(n_958),
.B1(n_984),
.B2(n_936),
.C1(n_924),
.C2(n_944),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_987),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_994),
.B(n_903),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_995),
.B(n_961),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_992),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_1001),
.B(n_983),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1004),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1022),
.B(n_1020),
.Y(n_1030)
);

AO21x2_ASAP7_75t_L g1031 ( 
.A1(n_1028),
.A2(n_1001),
.B(n_982),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_1011),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1029),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1029),
.Y(n_1034)
);

AO221x1_ASAP7_75t_L g1035 ( 
.A1(n_1023),
.A2(n_997),
.B1(n_1003),
.B2(n_962),
.C(n_960),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1022),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1011),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1017),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1015),
.B(n_1004),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1018),
.B(n_998),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1027),
.B(n_1005),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1019),
.Y(n_1043)
);

NAND2xp67_ASAP7_75t_L g1044 ( 
.A(n_1038),
.B(n_956),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1032),
.B(n_1012),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_1035),
.A2(n_1010),
.B1(n_1009),
.B2(n_1025),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1033),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1034),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1032),
.B(n_1012),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1031),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1040),
.B(n_1010),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1041),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1047),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1052),
.B(n_1030),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1048),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1045),
.B(n_1040),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1051),
.B(n_1036),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1049),
.Y(n_1058)
);

BUFx2_ASAP7_75t_SL g1059 ( 
.A(n_1058),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1053),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1056),
.B(n_1051),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1055),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1054),
.Y(n_1063)
);

OAI31xp33_ASAP7_75t_SL g1064 ( 
.A1(n_1057),
.A2(n_1046),
.A3(n_1028),
.B(n_1050),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1053),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_1056),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1058),
.B(n_1046),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_1014),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1061),
.B(n_1014),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1063),
.B(n_1037),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1061),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1060),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_1064),
.B(n_1050),
.C(n_1039),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1067),
.B(n_1031),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_1068),
.C(n_1066),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_1059),
.Y(n_1078)
);

AOI221x1_ASAP7_75t_L g1079 ( 
.A1(n_1071),
.A2(n_1065),
.B1(n_1062),
.B2(n_1068),
.C(n_1041),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1071),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1076),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_SL g1082 ( 
.A(n_1074),
.B(n_983),
.C(n_1026),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1073),
.A2(n_1043),
.B1(n_937),
.B2(n_949),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1080),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1079),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1081),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1078),
.B(n_1069),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1077),
.B(n_1069),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

XNOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1085),
.B(n_1072),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1085),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1087),
.B(n_1082),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1086),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1084),
.B(n_974),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1091),
.A2(n_1083),
.B(n_985),
.C(n_1042),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1089),
.A2(n_870),
.B(n_877),
.C(n_790),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1090),
.A2(n_974),
.B1(n_767),
.B2(n_951),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1094),
.Y(n_1098)
);

OAI211xp5_ASAP7_75t_L g1099 ( 
.A1(n_1093),
.A2(n_889),
.B(n_997),
.C(n_790),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1094),
.B(n_1044),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1098),
.B(n_1092),
.C(n_934),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_977),
.B1(n_936),
.B2(n_924),
.Y(n_1102)
);

AOI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1095),
.A2(n_1024),
.B1(n_1019),
.B2(n_941),
.C1(n_947),
.C2(n_1000),
.Y(n_1103)
);

AOI211x1_ASAP7_75t_SL g1104 ( 
.A1(n_1099),
.A2(n_1024),
.B(n_1021),
.C(n_1016),
.Y(n_1104)
);

OAI211xp5_ASAP7_75t_L g1105 ( 
.A1(n_1097),
.A2(n_1021),
.B(n_1016),
.C(n_1003),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_1101),
.Y(n_1107)
);

OAI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1103),
.A2(n_1096),
.B1(n_943),
.B2(n_949),
.C(n_935),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1105),
.B(n_977),
.Y(n_1109)
);

XOR2x1_ASAP7_75t_L g1110 ( 
.A(n_1102),
.B(n_948),
.Y(n_1110)
);

OAI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1104),
.A2(n_935),
.B1(n_762),
.B2(n_948),
.C(n_918),
.Y(n_1111)
);

OAI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1101),
.A2(n_762),
.B(n_786),
.C(n_962),
.Y(n_1112)
);

OAI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1104),
.A2(n_786),
.B1(n_787),
.B2(n_761),
.C(n_759),
.Y(n_1113)
);

NOR3x1_ASAP7_75t_L g1114 ( 
.A(n_1106),
.B(n_928),
.C(n_856),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1107),
.A2(n_857),
.B(n_875),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1112),
.B(n_161),
.C(n_162),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1109),
.A2(n_896),
.B(n_844),
.C(n_846),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1110),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1108),
.A2(n_969),
.B1(n_884),
.B2(n_927),
.Y(n_1119)
);

OAI322xp33_ASAP7_75t_L g1120 ( 
.A1(n_1111),
.A2(n_947),
.A3(n_996),
.B1(n_990),
.B2(n_988),
.C1(n_789),
.C2(n_772),
.Y(n_1120)
);

OAI321xp33_ASAP7_75t_L g1121 ( 
.A1(n_1113),
.A2(n_759),
.A3(n_761),
.B1(n_787),
.B2(n_986),
.C(n_911),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1107),
.B(n_969),
.Y(n_1122)
);

OAI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1106),
.A2(n_928),
.B(n_972),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_SL g1124 ( 
.A(n_1118),
.B(n_769),
.C(n_772),
.Y(n_1124)
);

AOI211xp5_ASAP7_75t_L g1125 ( 
.A1(n_1120),
.A2(n_849),
.B(n_842),
.C(n_862),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_1122),
.B(n_163),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1114),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_972),
.B1(n_911),
.B2(n_946),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_1115),
.B(n_884),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1116),
.A2(n_946),
.B1(n_911),
.B2(n_789),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1119),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1117),
.Y(n_1132)
);

NAND4xp25_ASAP7_75t_L g1133 ( 
.A(n_1121),
.B(n_780),
.C(n_902),
.D(n_899),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_1118),
.Y(n_1134)
);

AND3x1_ASAP7_75t_L g1135 ( 
.A(n_1118),
.B(n_996),
.C(n_990),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1116),
.B(n_988),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1127),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1126),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1132),
.Y(n_1139)
);

NAND4xp25_ASAP7_75t_L g1140 ( 
.A(n_1134),
.B(n_780),
.C(n_165),
.D(n_166),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_1124),
.B(n_164),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1135),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1136),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1133),
.A2(n_931),
.B(n_911),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1129),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1137),
.A2(n_1131),
.B1(n_1130),
.B2(n_1125),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1138),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1139),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_SL g1149 ( 
.A1(n_1142),
.A2(n_1128),
.B1(n_761),
.B2(n_787),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1139),
.Y(n_1150)
);

XNOR2xp5_ASAP7_75t_L g1151 ( 
.A(n_1140),
.B(n_167),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1143),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

AND2x2_ASAP7_75t_SL g1154 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1147),
.B(n_1152),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1155),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_1156),
.B(n_1153),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1157),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1158),
.A2(n_1154),
.B1(n_1146),
.B2(n_1149),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1158),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1158),
.A2(n_1145),
.B1(n_1144),
.B2(n_1141),
.C(n_946),
.Y(n_1161)
);

AOI222xp33_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_946),
.B1(n_911),
.B2(n_172),
.C1(n_173),
.C2(n_174),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1159),
.A2(n_920),
.B(n_904),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1161),
.B(n_946),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_1160),
.A2(n_168),
.B1(n_171),
.B2(n_175),
.C1(n_176),
.C2(n_178),
.Y(n_1165)
);

OAI22x1_ASAP7_75t_L g1166 ( 
.A1(n_1164),
.A2(n_179),
.B1(n_181),
.B2(n_183),
.Y(n_1166)
);

AOI222xp33_ASAP7_75t_L g1167 ( 
.A1(n_1163),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.C1(n_188),
.C2(n_193),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1165),
.A2(n_1162),
.B1(n_931),
.B2(n_197),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1164),
.A2(n_927),
.B1(n_904),
.B2(n_920),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1168),
.A2(n_195),
.B(n_196),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1166),
.B(n_925),
.Y(n_1171)
);

AO221x1_ASAP7_75t_L g1172 ( 
.A1(n_1167),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.C(n_204),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1170),
.A2(n_1169),
.B1(n_205),
.B2(n_206),
.C(n_207),
.Y(n_1173)
);

AOI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1173),
.A2(n_1171),
.B(n_1172),
.C(n_209),
.Y(n_1174)
);


endmodule