module fake_netlist_6_2871_n_70 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_70);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_70;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_18;
wire n_21;
wire n_24;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_64;
wire n_30;
wire n_43;
wire n_19;
wire n_48;
wire n_47;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_40;
wire n_25;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_13),
.B1(n_9),
.B2(n_14),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

OAI22x1_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_4),
.B1(n_9),
.B2(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_10),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_1),
.A2(n_2),
.B1(n_16),
.B2(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_22),
.Y(n_32)
);

NAND3x1_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_31),
.C(n_28),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_35),
.C(n_34),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_27),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_18),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_25),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_56),
.Y(n_59)
);

AOI222xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_49),
.B1(n_54),
.B2(n_21),
.C1(n_50),
.C2(n_47),
.Y(n_60)
);

NOR4xp25_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_46),
.C(n_25),
.D(n_51),
.Y(n_61)
);

AND4x1_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_51),
.C(n_25),
.D(n_57),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_51),
.B(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_59),
.C(n_57),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_30),
.B1(n_24),
.B2(n_45),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_25),
.C(n_63),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_61),
.B(n_52),
.Y(n_68)
);

AOI221x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_30),
.B1(n_66),
.B2(n_52),
.C(n_25),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_52),
.Y(n_70)
);


endmodule