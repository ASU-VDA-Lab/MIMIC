module fake_netlist_1_793_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_25;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_8), .B(n_7), .Y(n_13) );
BUFx10_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
BUFx10_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_1), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g20 ( .A(n_13), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_19), .B(n_2), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_15), .B(n_4), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_SL g25 ( .A1(n_15), .A2(n_9), .B(n_7), .C(n_8), .Y(n_25) );
BUFx8_ASAP7_75t_SL g26 ( .A(n_24), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_23), .B(n_13), .Y(n_28) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_21), .B(n_18), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NOR3xp33_ASAP7_75t_L g31 ( .A(n_30), .B(n_20), .C(n_29), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_28), .B1(n_12), .B2(n_17), .C1(n_16), .C2(n_27), .Y(n_33) );
INVxp67_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
CKINVDCx16_ASAP7_75t_R g35 ( .A(n_33), .Y(n_35) );
A2O1A1Ixp33_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_25), .B(n_16), .C(n_14), .Y(n_36) );
OAI22x1_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_26), .B1(n_25), .B2(n_5), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
AOI22xp5_ASAP7_75t_SL g39 ( .A1(n_37), .A2(n_5), .B1(n_14), .B2(n_38), .Y(n_39) );
endmodule