module fake_jpeg_6373_n_65 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_62;
wire n_56;
wire n_31;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_48),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_17),
.B1(n_29),
.B2(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_18),
.B1(n_28),
.B2(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_19),
.B1(n_7),
.B2(n_8),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_20),
.B1(n_9),
.B2(n_10),
.Y(n_48)
);

CKINVDCx10_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2x1_ASAP7_75t_R g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

XNOR2x1_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_1),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_39),
.B2(n_31),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.CI(n_52),
.CON(n_60),
.SN(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_34),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_60),
.C(n_32),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_12),
.B(n_13),
.Y(n_63)
);

AOI211xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_22),
.B(n_24),
.C(n_26),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_27),
.Y(n_65)
);


endmodule