module fake_jpeg_15619_n_15 (n_3, n_2, n_1, n_0, n_4, n_15);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_15;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

CKINVDCx12_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_0),
.Y(n_9)
);

AO221x1_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.C(n_7),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g11 ( 
.A1(n_5),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_5),
.Y(n_14)
);

OAI31xp33_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_6),
.A3(n_12),
.B(n_13),
.Y(n_15)
);


endmodule