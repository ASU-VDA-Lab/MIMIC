module fake_jpeg_2906_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_6),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_9),
.B1(n_13),
.B2(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_11),
.B1(n_22),
.B2(n_28),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_11),
.B1(n_18),
.B2(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_18),
.B1(n_21),
.B2(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_45),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_32),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_40),
.B(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_37),
.C(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_31),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.C(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_44),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_42),
.C(n_47),
.Y(n_53)
);

AOI31xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_47),
.A3(n_49),
.B(n_45),
.Y(n_54)
);


endmodule