module fake_jpeg_27106_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_16),
.B1(n_21),
.B2(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_9),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_21),
.B1(n_15),
.B2(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_14),
.B(n_7),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_14),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_19),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_34)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

MAJx2_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_29),
.C(n_28),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_33),
.B1(n_19),
.B2(n_10),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_11),
.B1(n_3),
.B2(n_6),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_33),
.B(n_5),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_41),
.C(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_5),
.Y(n_47)
);


endmodule