module real_aes_18100_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g825 ( .A(n_0), .B(n_826), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_1), .A2(n_3), .B1(n_181), .B2(n_524), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_2), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_4), .A2(n_44), .B1(n_138), .B2(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_5), .A2(n_119), .B1(n_120), .B2(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_5), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_481), .B1(n_486), .B2(n_488), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_6), .A2(n_27), .B1(n_161), .B2(n_237), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_7), .A2(n_17), .B1(n_180), .B2(n_216), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_8), .A2(n_61), .B1(n_198), .B2(n_239), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_9), .A2(n_18), .B1(n_137), .B2(n_138), .Y(n_540) );
INVx1_ASAP7_75t_L g826 ( .A(n_10), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_11), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_12), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_13), .A2(n_20), .B1(n_197), .B2(n_200), .Y(n_196) );
OR2x2_ASAP7_75t_L g111 ( .A(n_14), .B(n_40), .Y(n_111) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_15), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_16), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_19), .A2(n_100), .B1(n_820), .B2(n_830), .Y(n_99) );
OAI22xp33_ASAP7_75t_L g118 ( .A1(n_21), .A2(n_119), .B1(n_120), .B2(n_467), .Y(n_118) );
INVx2_ASAP7_75t_L g467 ( .A(n_21), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_22), .A2(n_97), .B1(n_180), .B2(n_181), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_23), .A2(n_41), .B1(n_146), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_24), .B(n_141), .Y(n_140) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_25), .A2(n_58), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_26), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_28), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_29), .B(n_143), .Y(n_510) );
INVx4_ASAP7_75t_R g552 ( .A(n_30), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_31), .A2(n_48), .B1(n_166), .B2(n_167), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_32), .A2(n_54), .B1(n_167), .B2(n_180), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_33), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_34), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_35), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_36), .B(n_161), .Y(n_517) );
INVx1_ASAP7_75t_L g526 ( .A(n_37), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_SL g592 ( .A1(n_38), .A2(n_138), .B(n_142), .C(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_39), .A2(n_55), .B1(n_138), .B2(n_167), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_42), .A2(n_85), .B1(n_138), .B2(n_236), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_43), .A2(n_47), .B1(n_137), .B2(n_138), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_45), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_46), .A2(n_60), .B1(n_180), .B2(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g514 ( .A(n_49), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_50), .B(n_138), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_51), .Y(n_573) );
INVx2_ASAP7_75t_L g115 ( .A(n_52), .Y(n_115) );
INVx1_ASAP7_75t_L g109 ( .A(n_53), .Y(n_109) );
BUFx3_ASAP7_75t_L g479 ( .A(n_53), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_56), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_57), .A2(n_86), .B1(n_138), .B2(n_167), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_59), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_62), .A2(n_74), .B1(n_166), .B2(n_184), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_63), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_64), .A2(n_76), .B1(n_137), .B2(n_138), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_65), .A2(n_95), .B1(n_180), .B2(n_200), .Y(n_226) );
INVx1_ASAP7_75t_L g133 ( .A(n_66), .Y(n_133) );
AND2x4_ASAP7_75t_L g152 ( .A(n_67), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_68), .A2(n_88), .B1(n_166), .B2(n_167), .Y(n_522) );
AO22x1_ASAP7_75t_L g531 ( .A1(n_69), .A2(n_75), .B1(n_213), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g153 ( .A(n_70), .Y(n_153) );
AND2x2_ASAP7_75t_L g595 ( .A(n_71), .B(n_155), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_72), .B(n_239), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_73), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_77), .B(n_161), .Y(n_574) );
INVx2_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_79), .B(n_155), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_80), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_81), .A2(n_96), .B1(n_167), .B2(n_239), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_82), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_83), .B(n_188), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_84), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_87), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_89), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_90), .B(n_155), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g473 ( .A(n_91), .Y(n_473) );
NAND2xp33_ASAP7_75t_L g148 ( .A(n_92), .B(n_141), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_93), .A2(n_203), .B(n_239), .C(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g554 ( .A(n_94), .B(n_555), .Y(n_554) );
NAND2xp33_ASAP7_75t_L g578 ( .A(n_98), .B(n_147), .Y(n_578) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_112), .Y(n_100) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_101), .A2(n_117), .B(n_118), .Y(n_116) );
NOR2x1_ASAP7_75t_R g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx4_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx8_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_106), .Y(n_117) );
AND2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_109), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_110), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1_ASAP7_75t_L g819 ( .A(n_111), .B(n_479), .Y(n_819) );
BUFx2_ASAP7_75t_L g829 ( .A(n_111), .Y(n_829) );
OAI21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_468), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g476 ( .A(n_115), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_115), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_411), .Y(n_121) );
NOR3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_329), .C(n_366), .Y(n_122) );
NAND4xp75_ASAP7_75t_L g123 ( .A(n_124), .B(n_249), .C(n_283), .D(n_313), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI32xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_171), .A3(n_221), .B1(n_230), .B2(n_244), .Y(n_125) );
OR2x2_ASAP7_75t_L g230 ( .A(n_126), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_127), .A2(n_441), .B(n_443), .Y(n_440) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_156), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_128), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g312 ( .A(n_128), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g407 ( .A(n_128), .B(n_223), .Y(n_407) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx2_ASAP7_75t_L g256 ( .A(n_129), .Y(n_256) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_129) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_289) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g155 ( .A(n_131), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_131), .B(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g218 ( .A(n_131), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_131), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_131), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g518 ( .A(n_131), .B(n_501), .Y(n_518) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_144), .B(n_150), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_140), .C(n_142), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g572 ( .A1(n_137), .A2(n_573), .B(n_574), .C(n_575), .Y(n_572) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_139), .Y(n_141) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
INVx2_ASAP7_75t_L g237 ( .A(n_139), .Y(n_237) );
INVx1_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
INVx3_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_141), .Y(n_532) );
INVx6_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_142), .A2(n_531), .B(n_533), .C(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_142), .A2(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_142), .B(n_531), .Y(n_604) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
INVx1_ASAP7_75t_L g513 ( .A(n_143), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_149), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_147), .A2(n_217), .B1(n_552), .B2(n_553), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_149), .A2(n_160), .B1(n_162), .B2(n_165), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_162), .B1(n_179), .B2(n_183), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_196), .B1(n_201), .B2(n_202), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_149), .A2(n_162), .B1(n_212), .B2(n_215), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_149), .A2(n_202), .B1(n_226), .B2(n_227), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_149), .A2(n_235), .B1(n_238), .B2(n_240), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_149), .A2(n_162), .B1(n_274), .B2(n_275), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_149), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_149), .A2(n_240), .B1(n_522), .B2(n_523), .Y(n_521) );
OAI22x1_ASAP7_75t_L g539 ( .A1(n_149), .A2(n_240), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_SL g241 ( .A(n_151), .Y(n_241) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx10_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx10_ASAP7_75t_L g501 ( .A(n_152), .Y(n_501) );
INVx1_ASAP7_75t_L g537 ( .A(n_152), .Y(n_537) );
INVx2_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_155), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g280 ( .A(n_156), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_156), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_157), .Y(n_267) );
INVx1_ASAP7_75t_L g311 ( .A(n_157), .Y(n_311) );
AND2x2_ASAP7_75t_L g355 ( .A(n_157), .B(n_289), .Y(n_355) );
OR2x2_ASAP7_75t_L g409 ( .A(n_157), .B(n_233), .Y(n_409) );
AO31x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .A3(n_168), .B(n_169), .Y(n_157) );
INVx2_ASAP7_75t_L g177 ( .A(n_158), .Y(n_177) );
AO31x2_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_195), .A3(n_204), .B(n_206), .Y(n_194) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_211), .A3(n_218), .B(n_219), .Y(n_210) );
AO31x2_ASAP7_75t_L g538 ( .A1(n_158), .A2(n_191), .A3(n_539), .B(n_542), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_161), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g500 ( .A(n_163), .Y(n_500) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g576 ( .A(n_164), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_167), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g524 ( .A(n_167), .Y(n_524) );
AO31x2_ASAP7_75t_L g496 ( .A1(n_168), .A2(n_497), .A3(n_501), .B(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_172), .A2(n_335), .B1(n_427), .B2(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_192), .Y(n_172) );
INVx4_ASAP7_75t_L g252 ( .A(n_173), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_173), .A2(n_232), .B1(n_264), .B2(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g269 ( .A(n_173), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g388 ( .A(n_173), .B(n_287), .Y(n_388) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g308 ( .A(n_174), .B(n_193), .Y(n_308) );
AND2x2_ASAP7_75t_L g399 ( .A(n_174), .B(n_271), .Y(n_399) );
AND2x2_ASAP7_75t_L g454 ( .A(n_174), .B(n_210), .Y(n_454) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
AND2x4_ASAP7_75t_L g375 ( .A(n_175), .B(n_271), .Y(n_375) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .A3(n_185), .B(n_189), .Y(n_175) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_176), .A2(n_204), .A3(n_225), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_177), .A2(n_547), .B(n_550), .Y(n_546) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_182), .B(n_590), .Y(n_589) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_185), .A2(n_241), .A3(n_273), .B(n_276), .Y(n_272) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_185), .A2(n_546), .B(n_554), .Y(n_545) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_SL g206 ( .A(n_187), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_187), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g191 ( .A(n_188), .Y(n_191) );
INVx2_ASAP7_75t_L g205 ( .A(n_188), .Y(n_205) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_188), .A2(n_535), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_191), .B(n_277), .Y(n_276) );
NAND2x1_ASAP7_75t_L g251 ( .A(n_192), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_192), .B(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
INVx2_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_193), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_193), .B(n_296), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_193), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g384 ( .A(n_193), .Y(n_384) );
INVx4_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_194), .B(n_209), .Y(n_262) );
BUFx2_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
AND2x2_ASAP7_75t_L g349 ( .A(n_194), .B(n_210), .Y(n_349) );
AND2x2_ASAP7_75t_L g391 ( .A(n_194), .B(n_272), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_194), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_199), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_204), .A2(n_241), .A3(n_521), .B(n_525), .Y(n_520) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_204), .A2(n_585), .B(n_595), .Y(n_584) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_205), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_205), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_205), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g555 ( .A(n_205), .Y(n_555) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_210), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g302 ( .A(n_210), .B(n_272), .Y(n_302) );
INVx1_ASAP7_75t_L g325 ( .A(n_210), .Y(n_325) );
INVx2_ASAP7_75t_L g345 ( .A(n_210), .Y(n_345) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_210), .Y(n_390) );
OAI21xp33_ASAP7_75t_SL g509 ( .A1(n_213), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AO31x2_ASAP7_75t_L g233 ( .A1(n_218), .A2(n_234), .A3(n_241), .B(n_242), .Y(n_233) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g309 ( .A(n_222), .B(n_310), .Y(n_309) );
NOR2x1p5_ASAP7_75t_L g415 ( .A(n_222), .B(n_409), .Y(n_415) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g232 ( .A(n_223), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_223), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_223), .B(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g257 ( .A(n_224), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g315 ( .A(n_224), .B(n_233), .Y(n_315) );
BUFx2_ASAP7_75t_L g428 ( .A(n_224), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_230), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g466 ( .A(n_230), .Y(n_466) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g402 ( .A(n_232), .Y(n_402) );
AND2x4_ASAP7_75t_L g425 ( .A(n_232), .B(n_355), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_232), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
BUFx2_ASAP7_75t_L g282 ( .A(n_233), .Y(n_282) );
INVx1_ASAP7_75t_L g338 ( .A(n_233), .Y(n_338) );
OR2x2_ASAP7_75t_L g460 ( .A(n_233), .B(n_317), .Y(n_460) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_237), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_240), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_247), .Y(n_323) );
INVx1_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
OR2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_297), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B(n_259), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_254), .A2(n_348), .B1(n_350), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OR2x2_ASAP7_75t_L g393 ( .A(n_256), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_256), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_256), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g376 ( .A(n_257), .B(n_355), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B1(n_269), .B2(n_278), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g328 ( .A(n_262), .Y(n_328) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g286 ( .A(n_265), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g354 ( .A(n_265), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g363 ( .A(n_265), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_265), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g351 ( .A(n_268), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g365 ( .A(n_268), .Y(n_365) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g297 ( .A(n_272), .Y(n_297) );
AND2x4_ASAP7_75t_L g344 ( .A(n_272), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_272), .Y(n_360) );
INVx1_ASAP7_75t_L g424 ( .A(n_272), .Y(n_424) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x4_ASAP7_75t_L g316 ( .A(n_280), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g333 ( .A(n_280), .Y(n_333) );
INVx1_ASAP7_75t_L g291 ( .A(n_282), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_292), .B1(n_303), .B2(n_309), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_288), .Y(n_341) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_298), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_294), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g446 ( .A(n_295), .Y(n_446) );
INVx1_ASAP7_75t_L g465 ( .A(n_295), .Y(n_465) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_299), .B(n_365), .Y(n_442) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g458 ( .A(n_300), .Y(n_458) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
INVx2_ASAP7_75t_L g396 ( .A(n_304), .Y(n_396) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g385 ( .A(n_305), .Y(n_385) );
AND2x4_ASAP7_75t_L g387 ( .A(n_306), .B(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_310), .A2(n_456), .B1(n_459), .B2(n_461), .Y(n_455) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g380 ( .A(n_311), .Y(n_380) );
INVx1_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
AND2x4_ASAP7_75t_L g427 ( .A(n_312), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g435 ( .A(n_312), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_318), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_SL g378 ( .A(n_315), .Y(n_378) );
INVx2_ASAP7_75t_L g394 ( .A(n_315), .Y(n_394) );
INVx1_ASAP7_75t_L g421 ( .A(n_316), .Y(n_421) );
AND2x2_ASAP7_75t_L g452 ( .A(n_316), .B(n_363), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .C(n_326), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_323), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g364 ( .A(n_324), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_324), .B(n_399), .Y(n_432) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_327), .B(n_391), .Y(n_417) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_346), .C(n_356), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B(n_342), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g450 ( .A(n_333), .Y(n_450) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g386 ( .A1(n_337), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_392), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_337), .B(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_344), .B(n_365), .Y(n_405) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_349), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g410 ( .A(n_349), .B(n_359), .Y(n_410) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g438 ( .A(n_352), .Y(n_438) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_354), .A2(n_357), .B1(n_361), .B2(n_364), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_355), .B(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_357), .A2(n_415), .B1(n_452), .B2(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g453 ( .A(n_359), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_361), .A2(n_404), .B1(n_406), .B2(n_410), .Y(n_403) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g445 ( .A(n_365), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_386), .C(n_395), .D(n_403), .Y(n_366) );
O2A1O1Ixp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_373), .B(n_376), .C(n_377), .Y(n_367) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g431 ( .A(n_375), .B(n_390), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_375), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_382), .A2(n_420), .B1(n_422), .B2(n_425), .Y(n_419) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_387), .A2(n_392), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_400), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_R g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_410), .A2(n_427), .B1(n_464), .B2(n_466), .Y(n_463) );
NOR3x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_433), .C(n_447), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_426), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
INVx1_ASAP7_75t_L g436 ( .A(n_428), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_430), .A2(n_434), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g447 ( .A(n_448), .B(n_451), .C(n_455), .D(n_463), .Y(n_447) );
AND2x2_ASAP7_75t_L g461 ( .A(n_454), .B(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI221x1_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_480), .B1(n_482), .B2(n_485), .C(n_811), .Y(n_468) );
NOR2xp67_ASAP7_75t_SL g469 ( .A(n_470), .B(n_474), .Y(n_469) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g818 ( .A(n_472), .B(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g484 ( .A(n_473), .Y(n_484) );
NOR2x1_ASAP7_75t_R g482 ( .A(n_474), .B(n_483), .Y(n_482) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_SL g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g823 ( .A(n_484), .B(n_824), .C(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_688), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_636), .Y(n_489) );
OAI211xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_527), .B(n_556), .C(n_621), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_493), .A2(n_557), .B(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
INVx2_ASAP7_75t_L g617 ( .A(n_494), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_494), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g728 ( .A(n_495), .B(n_506), .Y(n_728) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g596 ( .A(n_496), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_496), .B(n_520), .Y(n_633) );
AND2x2_ASAP7_75t_L g666 ( .A(n_496), .B(n_583), .Y(n_666) );
OR2x2_ASAP7_75t_L g671 ( .A(n_496), .B(n_520), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_500), .A2(n_516), .B(n_517), .Y(n_515) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_500), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g581 ( .A(n_501), .Y(n_581) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g810 ( .A(n_505), .Y(n_810) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_519), .Y(n_505) );
AND2x2_ASAP7_75t_L g611 ( .A(n_506), .B(n_520), .Y(n_611) );
INVx3_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
NAND2x1p5_ASAP7_75t_SL g651 ( .A(n_506), .B(n_635), .Y(n_651) );
INVx1_ASAP7_75t_L g669 ( .A(n_506), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_506), .B(n_614), .Y(n_694) );
BUFx2_ASAP7_75t_L g780 ( .A(n_506), .Y(n_780) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_515), .B(n_518), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_513), .Y(n_591) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
INVx1_ASAP7_75t_L g620 ( .A(n_520), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_520), .B(n_596), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_520), .B(n_583), .Y(n_729) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_544), .Y(n_527) );
INVx1_ASAP7_75t_L g787 ( .A(n_528), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
OR2x2_ASAP7_75t_L g559 ( .A(n_529), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g624 ( .A(n_529), .Y(n_624) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g603 ( .A(n_533), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_536), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_537), .A2(n_586), .B(n_592), .Y(n_585) );
INVx2_ASAP7_75t_L g560 ( .A(n_538), .Y(n_560) );
OR2x2_ASAP7_75t_L g625 ( .A(n_538), .B(n_545), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_538), .B(n_545), .Y(n_630) );
INVx2_ASAP7_75t_L g675 ( .A(n_538), .Y(n_675) );
AND2x2_ASAP7_75t_L g716 ( .A(n_538), .B(n_569), .Y(n_716) );
AND2x2_ASAP7_75t_L g750 ( .A(n_538), .B(n_647), .Y(n_750) );
INVx1_ASAP7_75t_L g561 ( .A(n_544), .Y(n_561) );
INVx1_ASAP7_75t_L g680 ( .A(n_544), .Y(n_680) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g600 ( .A(n_545), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g641 ( .A(n_545), .B(n_602), .Y(n_641) );
INVx2_ASAP7_75t_L g647 ( .A(n_545), .Y(n_647) );
AND2x2_ASAP7_75t_L g702 ( .A(n_545), .B(n_569), .Y(n_702) );
AND2x2_ASAP7_75t_L g759 ( .A(n_545), .B(n_568), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_562), .B1(n_597), .B2(n_608), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
NAND3xp33_ASAP7_75t_SL g737 ( .A(n_559), .B(n_738), .C(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g656 ( .A(n_560), .Y(n_656) );
AND2x2_ASAP7_75t_L g706 ( .A(n_560), .B(n_568), .Y(n_706) );
INVx1_ASAP7_75t_L g806 ( .A(n_561), .Y(n_806) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_563), .B(n_761), .Y(n_797) );
BUFx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g652 ( .A(n_564), .Y(n_652) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_582), .Y(n_566) );
INVx1_ASAP7_75t_L g640 ( .A(n_567), .Y(n_640) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g720 ( .A(n_568), .B(n_601), .Y(n_720) );
AND2x2_ASAP7_75t_L g739 ( .A(n_568), .B(n_646), .Y(n_739) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g607 ( .A(n_569), .Y(n_607) );
BUFx3_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g674 ( .A(n_569), .B(n_675), .Y(n_674) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B(n_580), .Y(n_571) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g767 ( .A(n_582), .Y(n_767) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_596), .Y(n_582) );
INVx2_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_591), .Y(n_586) );
INVx1_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_599), .B(n_606), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g654 ( .A(n_600), .B(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g784 ( .A(n_600), .Y(n_784) );
INVx1_ASAP7_75t_L g629 ( .A(n_601), .Y(n_629) );
AND2x2_ASAP7_75t_L g709 ( .A(n_601), .B(n_647), .Y(n_709) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g646 ( .A(n_602), .B(n_647), .Y(n_646) );
AOI21x1_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_607), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g742 ( .A(n_607), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_616), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_609), .A2(n_650), .B1(n_653), .B2(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_610), .A2(n_630), .B1(n_662), .B2(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
BUFx2_ASAP7_75t_SL g648 ( .A(n_611), .Y(n_648) );
AND2x4_ASAP7_75t_L g766 ( .A(n_611), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g775 ( .A(n_611), .Y(n_775) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g687 ( .A(n_613), .Y(n_687) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_614), .B(n_619), .Y(n_745) );
INVxp67_ASAP7_75t_L g774 ( .A(n_614), .Y(n_774) );
AND2x2_ASAP7_75t_L g779 ( .A(n_614), .B(n_645), .Y(n_779) );
OR2x2_ASAP7_75t_L g761 ( .A(n_615), .B(n_635), .Y(n_761) );
INVx1_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_617), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g681 ( .A(n_618), .B(n_666), .Y(n_681) );
AND2x4_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_619), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g665 ( .A(n_619), .Y(n_665) );
OR2x2_ASAP7_75t_L g760 ( .A(n_619), .B(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_626), .B(n_631), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g684 ( .A(n_623), .Y(n_684) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g678 ( .A(n_624), .B(n_675), .Y(n_678) );
INVx2_ASAP7_75t_L g802 ( .A(n_624), .Y(n_802) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND2x2_ASAP7_75t_L g731 ( .A(n_628), .B(n_674), .Y(n_731) );
AND2x2_ASAP7_75t_L g756 ( .A(n_628), .B(n_702), .Y(n_756) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g659 ( .A(n_629), .Y(n_659) );
AND2x2_ASAP7_75t_L g686 ( .A(n_630), .B(n_640), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_630), .B(n_685), .Y(n_698) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g783 ( .A(n_633), .Y(n_783) );
OR2x2_ASAP7_75t_L g799 ( .A(n_633), .B(n_694), .Y(n_799) );
INVx1_ASAP7_75t_L g723 ( .A(n_635), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_660), .C(n_682), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_642), .B1(n_643), .B2(n_648), .C(n_649), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g662 ( .A(n_641), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_641), .B(n_706), .Y(n_790) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_L g685 ( .A(n_645), .Y(n_685) );
AND3x1_ASAP7_75t_L g781 ( .A(n_645), .B(n_782), .C(n_783), .Y(n_781) );
AND2x2_ASAP7_75t_L g768 ( .A(n_646), .B(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g778 ( .A(n_646), .Y(n_778) );
INVxp67_ASAP7_75t_L g792 ( .A(n_648), .Y(n_792) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OR2x2_ASAP7_75t_L g747 ( .A(n_651), .B(n_671), .Y(n_747) );
INVx2_ASAP7_75t_L g782 ( .A(n_651), .Y(n_782) );
INVx1_ASAP7_75t_L g700 ( .A(n_652), .Y(n_700) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_654), .A2(n_702), .B(n_703), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_655), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g663 ( .A(n_656), .Y(n_663) );
OR2x2_ASAP7_75t_L g757 ( .A(n_656), .B(n_758), .Y(n_757) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g717 ( .A(n_659), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_659), .B(n_716), .Y(n_796) );
AND3x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_667), .C(n_672), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
AND2x2_ASAP7_75t_L g711 ( .A(n_663), .B(n_702), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_664), .A2(n_731), .B1(n_732), .B2(n_734), .Y(n_730) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI321xp33_ASAP7_75t_L g753 ( .A1(n_665), .A2(n_754), .A3(n_755), .B1(n_757), .B2(n_760), .C(n_762), .Y(n_753) );
AND2x2_ASAP7_75t_L g805 ( .A(n_665), .B(n_670), .Y(n_805) );
AND2x2_ASAP7_75t_L g703 ( .A(n_666), .B(n_669), .Y(n_703) );
INVx2_ASAP7_75t_L g712 ( .A(n_668), .Y(n_712) );
AND2x2_ASAP7_75t_L g721 ( .A(n_668), .B(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g733 ( .A(n_671), .B(n_723), .Y(n_733) );
INVx2_ASAP7_75t_L g765 ( .A(n_671), .Y(n_765) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_681), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g769 ( .A(n_675), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_678), .B(n_685), .Y(n_695) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_686), .B(n_687), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_685), .B(n_709), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_685), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g786 ( .A(n_685), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g754 ( .A(n_687), .Y(n_754) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_689), .B(n_751), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_713), .C(n_736), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_704), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B1(n_696), .B2(n_699), .C(n_701), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OR2x2_ASAP7_75t_L g744 ( .A(n_693), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_710), .B(n_712), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g741 ( .A(n_709), .B(n_742), .Y(n_741) );
OAI21xp33_ASAP7_75t_SL g724 ( .A1(n_710), .A2(n_725), .B(n_730), .Y(n_724) );
INVx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B(n_721), .C(n_724), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_715), .B(n_790), .Y(n_789) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_723), .B(n_765), .Y(n_764) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_726), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_743), .B1(n_746), .B2(n_748), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_745), .Y(n_808) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_788), .C(n_803), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_770), .Y(n_752) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
OAI21xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .B(n_768), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_776), .C(n_785), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AOI32xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .A3(n_780), .B1(n_781), .B2(n_784), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g804 ( .A(n_779), .B(n_805), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_791), .B(n_793), .Y(n_788) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI22x1_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B1(n_798), .B2(n_800), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI21xp33_ASAP7_75t_L g807 ( .A1(n_796), .A2(n_808), .B(n_809), .Y(n_807) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_806), .B(n_807), .Y(n_803) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx10_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx4_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx6f_ASAP7_75t_SL g831 ( .A(n_822), .Y(n_831) );
AND2x2_ASAP7_75t_SL g822 ( .A(n_823), .B(n_828), .Y(n_822) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
INVx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
endmodule