module fake_jpeg_3343_n_352 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_49),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_5),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_56),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_59),
.B(n_84),
.Y(n_124)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_6),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_67),
.Y(n_137)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_74),
.Y(n_139)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_7),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_7),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_7),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_8),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_87),
.B(n_90),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_10),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_91),
.B(n_96),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_33),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_11),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_61),
.A2(n_32),
.B1(n_41),
.B2(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_181)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_18),
.B1(n_40),
.B2(n_35),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_32),
.B1(n_41),
.B2(n_18),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_93),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_150),
.B1(n_51),
.B2(n_98),
.Y(n_160)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_63),
.A2(n_31),
.B1(n_38),
.B2(n_48),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_86),
.B1(n_76),
.B2(n_56),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_79),
.A2(n_31),
.B1(n_45),
.B2(n_47),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_158),
.B(n_165),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_102),
.B1(n_144),
.B2(n_112),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_56),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_73),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_168),
.C(n_173),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_47),
.B(n_48),
.C(n_60),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_166),
.B(n_180),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_75),
.C(n_55),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_144),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_57),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_187),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_101),
.A2(n_95),
.B(n_99),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_196),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_70),
.C(n_94),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_195),
.C(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_119),
.B(n_14),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_183),
.B(n_189),
.Y(n_221)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_120),
.B(n_11),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_13),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_13),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_13),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_115),
.B(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_105),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_162),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_106),
.Y(n_198)
);

NAND2x1_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_179),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_134),
.B(n_132),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_148),
.B(n_111),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_171),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

OR2x2_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_165),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_205),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_103),
.B1(n_107),
.B2(n_114),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_147),
.B1(n_138),
.B2(n_156),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_104),
.B1(n_131),
.B2(n_123),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_169),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_145),
.C(n_117),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_167),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_230),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_109),
.B1(n_173),
.B2(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_168),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_163),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_252),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_234),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_233),
.Y(n_258)
);

AOI22x1_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_174),
.B1(n_171),
.B2(n_175),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_255),
.B1(n_236),
.B2(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_195),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_254),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_184),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_178),
.Y(n_241)
);

OAI22x1_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_182),
.B1(n_169),
.B2(n_163),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_212),
.B1(n_213),
.B2(n_211),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_159),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_248),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_182),
.B1(n_167),
.B2(n_177),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_186),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_253),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_177),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_201),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_221),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_250),
.B(n_253),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_261),
.B(n_227),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_204),
.B(n_229),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_264),
.B1(n_267),
.B2(n_276),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_200),
.B1(n_224),
.B2(n_223),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_200),
.B1(n_226),
.B2(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_271),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_216),
.C(n_203),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_243),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_229),
.B1(n_218),
.B2(n_226),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_214),
.B1(n_219),
.B2(n_225),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_236),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_279),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_252),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_278),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_239),
.B1(n_242),
.B2(n_248),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_282),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_247),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_239),
.B1(n_244),
.B2(n_248),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_240),
.C(n_241),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_270),
.C(n_284),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_249),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_214),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_266),
.C(n_267),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_219),
.B(n_225),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_260),
.C(n_266),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_264),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_259),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_270),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_283),
.B(n_270),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_289),
.B1(n_281),
.B2(n_290),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_314),
.Y(n_321)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_298),
.A2(n_295),
.B1(n_300),
.B2(n_306),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_277),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_316),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_268),
.B1(n_288),
.B2(n_280),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_304),
.Y(n_320)
);

BUFx12f_ASAP7_75t_SL g326 ( 
.A(n_320),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_303),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_330),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_311),
.C(n_317),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_332),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_315),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_334),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_305),
.C(n_293),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_327),
.B1(n_318),
.B2(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_323),
.B1(n_322),
.B2(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_305),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_336),
.A2(n_338),
.B(n_339),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_340),
.B(n_335),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_341),
.B(n_342),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_282),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_343),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_346),
.A2(n_347),
.B(n_326),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_307),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_302),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_291),
.B(n_272),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_291),
.A3(n_269),
.B1(n_271),
.B2(n_273),
.C1(n_282),
.C2(n_304),
.Y(n_351)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_280),
.B(n_322),
.Y(n_352)
);


endmodule