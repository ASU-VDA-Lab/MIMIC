module fake_jpeg_29552_n_89 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_4),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_41),
.B1(n_34),
.B2(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_36),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_54),
.B1(n_7),
.B2(n_8),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_34),
.B(n_37),
.C(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_32),
.B1(n_38),
.B2(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_49),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_10),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_17),
.B(n_18),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_12),
.C(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_64),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_71),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_20),
.C(n_22),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_23),
.C(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_78),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_78),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_82),
.A3(n_83),
.B1(n_76),
.B2(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);


endmodule