module fake_jpeg_2384_n_143 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_5),
.Y(n_40)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_14),
.B1(n_19),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_48),
.B1(n_54),
.B2(n_20),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_14),
.B1(n_19),
.B2(n_25),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_27),
.B1(n_20),
.B2(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_15),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_63),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_29),
.B(n_22),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_69),
.B(n_74),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_35),
.C(n_23),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_50),
.C(n_69),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_29),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_49),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_23),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_0),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_28),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_56),
.B1(n_52),
.B2(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_65),
.B1(n_60),
.B2(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_68),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_42),
.A3(n_44),
.B1(n_41),
.B2(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_57),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_89),
.C(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_105),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_88),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_74),
.B(n_65),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_106),
.C(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_11),
.C(n_13),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_62),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_62),
.C(n_57),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_112),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_113),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_90),
.B1(n_80),
.B2(n_85),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_80),
.C(n_84),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_116),
.C(n_28),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_106),
.C(n_102),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_120),
.C(n_125),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_119),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_109),
.C(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_0),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_135),
.B(n_127),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_139),
.C(n_2),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_127),
.B(n_1),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_138),
.B(n_2),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_0),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_141),
.B1(n_139),
.B2(n_2),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_4),
.C(n_140),
.Y(n_143)
);


endmodule