module fake_jpeg_826_n_102 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_29),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_26),
.B1(n_28),
.B2(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_54),
.B1(n_31),
.B2(n_2),
.Y(n_61)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_1),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_48),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_25),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_2),
.B(n_3),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_11),
.C(n_22),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_56),
.B1(n_54),
.B2(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_77),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_79),
.C(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_70),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_12),
.B1(n_21),
.B2(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_15),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_9),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

AOI31xp67_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_95),
.A3(n_89),
.B(n_80),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_88),
.C(n_72),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_93),
.B(n_90),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_91),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_10),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_75),
.Y(n_102)
);


endmodule