module fake_jpeg_9900_n_5 (n_0, n_1, n_5);

input n_0;
input n_1;

output n_5;

wire n_2;
wire n_3;
wire n_4;

INVx3_ASAP7_75t_L g2 ( 
.A(n_1),
.Y(n_2)
);

AND2x6_ASAP7_75t_L g3 ( 
.A(n_1),
.B(n_0),
.Y(n_3)
);

FAx1_ASAP7_75t_SL g4 ( 
.A(n_3),
.B(n_0),
.CI(n_2),
.CON(n_4),
.SN(n_4)
);

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_4),
.B(n_0),
.Y(n_5)
);


endmodule