module fake_netlist_6_94_n_1698 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1698);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1698;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g159 ( 
.A(n_126),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_24),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_34),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_32),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_30),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_54),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_72),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_4),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_35),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_91),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_57),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_41),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_90),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_19),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_41),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_55),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_66),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_106),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_50),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_158),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_33),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_93),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_42),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_71),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_20),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_113),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_60),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_86),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_50),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_38),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_43),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_36),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_110),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_69),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_57),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_80),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_125),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_100),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_92),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_145),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_19),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_56),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_146),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_47),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_124),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_3),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_123),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_28),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_16),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_112),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_122),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_107),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_131),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_49),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_27),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_52),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_51),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_35),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_39),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_101),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_150),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_138),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_49),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_129),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_98),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_36),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_82),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_88),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_76),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_114),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_38),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_12),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_149),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_89),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_153),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_119),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_28),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_276),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_195),
.B(n_0),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_190),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_193),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_207),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_244),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_198),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_208),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_172),
.B(n_1),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_169),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_209),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_169),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_169),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_214),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_296),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_172),
.B(n_1),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_305),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_215),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_169),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_217),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_310),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_178),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_220),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_258),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_226),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_169),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_227),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_231),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_238),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_196),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_249),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_196),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_173),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_250),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_228),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_251),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_196),
.B(n_3),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_252),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_253),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_166),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_196),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_196),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_166),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_260),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_262),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_259),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_167),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_196),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_266),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_189),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_167),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_191),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_242),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_173),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_242),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_242),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_242),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_242),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_258),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_242),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_177),
.B(n_6),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_173),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_200),
.B(n_6),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_258),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_258),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_268),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_388),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_317),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_277),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_388),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_191),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_258),
.Y(n_405)
);

CKINVDCx8_ASAP7_75t_R g406 ( 
.A(n_316),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_197),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_197),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_324),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_324),
.B(n_177),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_329),
.B(n_161),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_342),
.A2(n_315),
.B1(n_314),
.B2(n_313),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_334),
.B(n_161),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_182),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_348),
.B(n_352),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_348),
.B(n_175),
.Y(n_430)
);

INVx6_ASAP7_75t_L g431 ( 
.A(n_318),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_318),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_381),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_175),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_357),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_328),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_336),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_387),
.B(n_182),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_398),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_398),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_319),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_398),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_458),
.A2(n_390),
.B1(n_347),
.B2(n_353),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_396),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_320),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_225),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_396),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_375),
.Y(n_484)
);

INVx4_ASAP7_75t_SL g485 ( 
.A(n_431),
.Y(n_485)
);

INVx8_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_405),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_395),
.B(n_355),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_453),
.B(n_326),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_453),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_408),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_327),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_405),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_395),
.B(n_355),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_426),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_395),
.B(n_378),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_396),
.A2(n_322),
.B1(n_344),
.B2(n_323),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

NOR2x1p5_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_228),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_406),
.Y(n_506)
);

INVx4_ASAP7_75t_SL g507 ( 
.A(n_431),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_459),
.A2(n_387),
.B1(n_200),
.B2(n_307),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_454),
.B(n_378),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_330),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_338),
.C(n_333),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_340),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_458),
.B(n_386),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

OAI21xp33_ASAP7_75t_SL g520 ( 
.A1(n_460),
.A2(n_206),
.B(n_201),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_392),
.B(n_369),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_457),
.B(n_386),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_459),
.A2(n_264),
.B1(n_292),
.B2(n_224),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_392),
.B(n_343),
.Y(n_524)
);

BUFx4f_ASAP7_75t_L g525 ( 
.A(n_457),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_457),
.B(n_345),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_460),
.B(n_349),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_432),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_409),
.B(n_350),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_194),
.C(n_186),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_185),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_409),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_457),
.B(n_351),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_457),
.B(n_358),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_423),
.A2(n_288),
.B1(n_270),
.B2(n_211),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_460),
.B(n_168),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_421),
.B(n_367),
.C(n_362),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_434),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_394),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_459),
.A2(n_254),
.B1(n_281),
.B2(n_289),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_392),
.B(n_343),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_415),
.B(n_356),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_434),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_398),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_394),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_415),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_394),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_435),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_459),
.B(n_361),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_401),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_407),
.B(n_159),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_402),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_L g569 ( 
.A1(n_407),
.A2(n_374),
.B(n_293),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_454),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_435),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_407),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_403),
.B(n_374),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_459),
.B(n_368),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_459),
.A2(n_212),
.B1(n_243),
.B2(n_248),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_459),
.A2(n_274),
.B1(n_291),
.B2(n_211),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_437),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_403),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_401),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_225),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_437),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_407),
.B(n_229),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_448),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_421),
.B(n_232),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_402),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_440),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_425),
.B(n_373),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_401),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_425),
.B(n_309),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_423),
.A2(n_341),
.B1(n_337),
.B2(n_335),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_440),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_401),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_402),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_401),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_430),
.B(n_325),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_450),
.B(n_221),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_438),
.A2(n_237),
.B1(n_308),
.B2(n_203),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_443),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_443),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_431),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_431),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_450),
.B(n_183),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_438),
.B(n_287),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_561),
.B(n_391),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_524),
.B(n_442),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_554),
.B(n_391),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_467),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_467),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_488),
.B(n_581),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_472),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_532),
.B(n_442),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_554),
.B(n_391),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_463),
.B(n_391),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_565),
.A2(n_461),
.B1(n_428),
.B2(n_417),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_468),
.B(n_443),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_524),
.B(n_406),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_491),
.B(n_406),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_492),
.Y(n_626)
);

INVx8_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_477),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_557),
.B(n_449),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_492),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_487),
.B(n_417),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_471),
.A2(n_239),
.B1(n_315),
.B2(n_314),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_481),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_464),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_497),
.B(n_417),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_496),
.B(n_406),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_572),
.B(n_428),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_481),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_572),
.B(n_462),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_525),
.B(n_410),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_575),
.A2(n_461),
.B1(n_428),
.B2(n_284),
.Y(n_641)
);

BUFx6f_ASAP7_75t_SL g642 ( 
.A(n_573),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_462),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_552),
.B(n_521),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_462),
.B(n_424),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_488),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_606),
.B(n_527),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_183),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_466),
.B(n_424),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_540),
.A2(n_461),
.B1(n_270),
.B2(n_424),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_516),
.B(n_424),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_492),
.A2(n_267),
.B1(n_163),
.B2(n_164),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_465),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_517),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_483),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_465),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_525),
.B(n_546),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_476),
.B(n_187),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_511),
.B(n_168),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_587),
.B(n_424),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_567),
.A2(n_444),
.B(n_452),
.C(n_447),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_534),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_534),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_555),
.B(n_187),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_585),
.A2(n_246),
.B1(n_313),
.B2(n_306),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_461),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_544),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_552),
.B(n_461),
.Y(n_670)
);

INVx6_ASAP7_75t_L g671 ( 
.A(n_505),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_522),
.A2(n_461),
.B1(n_279),
.B2(n_302),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_546),
.B(n_410),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_540),
.A2(n_225),
.B1(n_273),
.B2(n_257),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_511),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_506),
.B(n_221),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_439),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_489),
.B(n_439),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_489),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_490),
.B(n_439),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_490),
.B(n_439),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_493),
.B(n_448),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_499),
.B(n_448),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_501),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_546),
.B(n_448),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_607),
.A2(n_239),
.B1(n_246),
.B2(n_306),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_503),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_503),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_515),
.B(n_240),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_512),
.B(n_448),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_512),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_529),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_498),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_529),
.B(n_448),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_533),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_533),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_486),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_510),
.B(n_448),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_591),
.A2(n_302),
.B1(n_240),
.B2(n_241),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_521),
.B(n_259),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_500),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_484),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_573),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_484),
.B(n_259),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_573),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_502),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_540),
.A2(n_225),
.B1(n_210),
.B2(n_205),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_537),
.B(n_448),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_510),
.B(n_436),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_469),
.B(n_241),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_599),
.B(n_545),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_537),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_473),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_539),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_573),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_506),
.B(n_300),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_510),
.B(n_436),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_505),
.A2(n_300),
.B1(n_303),
.B2(n_312),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_539),
.Y(n_720)
);

NAND2x1_ASAP7_75t_L g721 ( 
.A(n_504),
.B(n_431),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_549),
.B(n_422),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_570),
.B(n_569),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_486),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_510),
.B(n_436),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_549),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_594),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_470),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_558),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_510),
.B(n_436),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_564),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_422),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_526),
.A2(n_312),
.B1(n_303),
.B2(n_162),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_532),
.B(n_192),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_571),
.Y(n_737)
);

AND2x6_ASAP7_75t_L g738 ( 
.A(n_571),
.B(n_574),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_574),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_576),
.B(n_422),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_518),
.B(n_204),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_576),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_536),
.A2(n_165),
.B1(n_255),
.B2(n_245),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_579),
.B(n_427),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_541),
.B(n_170),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_532),
.B(n_179),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_532),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_553),
.B(n_436),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_486),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_541),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_579),
.B(n_427),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_584),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_584),
.B(n_427),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_607),
.B(n_213),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_520),
.B(n_393),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_589),
.B(n_427),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_486),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_540),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_538),
.A2(n_180),
.B1(n_230),
.B2(n_202),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_553),
.B(n_436),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_589),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_590),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_474),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_600),
.B(n_216),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_647),
.B(n_601),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_721),
.A2(n_580),
.B(n_504),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_614),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_664),
.A2(n_595),
.B(n_603),
.C(n_602),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_757),
.A2(n_580),
.B(n_504),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_698),
.B(n_553),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_758),
.A2(n_478),
.B(n_583),
.C(n_531),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_664),
.A2(n_603),
.B(n_602),
.C(n_523),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_643),
.B(n_553),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_757),
.A2(n_604),
.B(n_580),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_670),
.B(n_631),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_611),
.A2(n_605),
.B(n_604),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_611),
.A2(n_605),
.B(n_604),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_698),
.B(n_553),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_703),
.B(n_480),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_613),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_620),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_674),
.A2(n_577),
.B1(n_551),
.B2(n_508),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_641),
.A2(n_578),
.B1(n_605),
.B2(n_586),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_609),
.B(n_171),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_712),
.A2(n_583),
.B(n_304),
.C(n_299),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_645),
.A2(n_586),
.B(n_519),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_618),
.A2(n_586),
.B(n_519),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_698),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_624),
.B(n_485),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_712),
.A2(n_528),
.B1(n_475),
.B2(n_588),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_625),
.A2(n_528),
.B1(n_475),
.B2(n_588),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_705),
.B(n_171),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_635),
.B(n_597),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_495),
.B(n_568),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_668),
.B(n_474),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_675),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_655),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_620),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_724),
.A2(n_495),
.B(n_568),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_625),
.B(n_636),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_758),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_724),
.A2(n_495),
.B(n_568),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_724),
.A2(n_495),
.B(n_568),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_648),
.A2(n_188),
.B(n_199),
.C(n_280),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_728),
.B(n_676),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_749),
.A2(n_657),
.B(n_608),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_632),
.B(n_639),
.C(n_637),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_684),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_648),
.B(n_479),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_749),
.B(n_507),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_658),
.B(n_479),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_658),
.A2(n_741),
.B(n_690),
.C(n_764),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_649),
.A2(n_482),
.B(n_494),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_617),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_646),
.B(n_218),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_620),
.B(n_507),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_673),
.A2(n_598),
.B(n_596),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_667),
.B(n_283),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_621),
.A2(n_285),
.B1(n_295),
.B2(n_297),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_612),
.B(n_482),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_692),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_694),
.B(n_219),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_741),
.A2(n_598),
.B(n_596),
.C(n_592),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_620),
.B(n_507),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_673),
.A2(n_592),
.B(n_582),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_690),
.A2(n_582),
.B(n_566),
.C(n_563),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_701),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_692),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_615),
.B(n_494),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_651),
.A2(n_509),
.B(n_514),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_660),
.A2(n_661),
.B(n_682),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_702),
.B(n_548),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_739),
.B(n_507),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_667),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_640),
.A2(n_566),
.B(n_563),
.Y(n_838)
);

BUFx12f_ASAP7_75t_L g839 ( 
.A(n_617),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_683),
.A2(n_547),
.B(n_514),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_627),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_726),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_685),
.A2(n_562),
.B(n_560),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_685),
.A2(n_559),
.B(n_550),
.Y(n_844)
);

INVx5_ASAP7_75t_L g845 ( 
.A(n_738),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_666),
.A2(n_632),
.B(n_616),
.C(n_628),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_737),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_623),
.B(n_509),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_633),
.B(n_638),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_626),
.B(n_548),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_737),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_739),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_627),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_762),
.B(n_535),
.Y(n_854)
);

AO21x1_ASAP7_75t_L g855 ( 
.A1(n_743),
.A2(n_759),
.B(n_652),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_762),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_677),
.B(n_535),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_619),
.A2(n_416),
.B(n_542),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_717),
.B(n_221),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_747),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_622),
.B(n_542),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_691),
.A2(n_547),
.B(n_452),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_627),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_654),
.A2(n_452),
.B1(n_441),
.B2(n_447),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_764),
.B(n_719),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_678),
.A2(n_416),
.B(n_402),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_727),
.B(n_671),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_680),
.A2(n_416),
.B(n_402),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_745),
.B(n_247),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_659),
.B(n_706),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_679),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_716),
.B(n_222),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_695),
.A2(n_445),
.B(n_444),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_629),
.A2(n_445),
.B(n_444),
.C(n_441),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_642),
.B(n_176),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_681),
.A2(n_411),
.B(n_418),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_662),
.A2(n_411),
.B(n_418),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_754),
.B(n_176),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_699),
.A2(n_411),
.B(n_418),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_709),
.A2(n_445),
.B(n_414),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_738),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_663),
.B(n_436),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_723),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_710),
.A2(n_411),
.B(n_413),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_617),
.Y(n_885)
);

O2A1O1Ixp5_ASAP7_75t_L g886 ( 
.A1(n_687),
.A2(n_393),
.B(n_397),
.C(n_400),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_688),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_710),
.A2(n_411),
.B(n_413),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_750),
.B(n_223),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_750),
.B(n_233),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_665),
.B(n_436),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_718),
.A2(n_411),
.B(n_413),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_738),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_736),
.B(n_181),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_738),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_718),
.A2(n_414),
.B(n_419),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_689),
.B(n_693),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_696),
.B(n_436),
.Y(n_898)
);

NOR2x1_ASAP7_75t_R g899 ( 
.A(n_671),
.B(n_181),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_745),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_722),
.A2(n_419),
.B(n_414),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_697),
.B(n_436),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_755),
.A2(n_393),
.B(n_397),
.C(n_400),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_713),
.B(n_446),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_725),
.A2(n_411),
.B(n_419),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_626),
.B(n_247),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_746),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_715),
.B(n_446),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_711),
.B(n_286),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_725),
.A2(n_411),
.B(n_431),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_738),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_720),
.B(n_446),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_669),
.B(n_446),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_671),
.A2(n_630),
.B1(n_729),
.B2(n_752),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_732),
.A2(n_411),
.B(n_446),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_630),
.A2(n_272),
.B1(n_235),
.B2(n_236),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_731),
.B1(n_742),
.B2(n_733),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_761),
.B(n_451),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_610),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_672),
.B(n_247),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_SL g921 ( 
.A1(n_748),
.A2(n_404),
.B(n_247),
.C(n_10),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_734),
.A2(n_404),
.B(n_234),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_760),
.A2(n_451),
.B(n_446),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_740),
.A2(n_404),
.B(n_446),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_746),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_746),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_700),
.B(n_247),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_744),
.A2(n_451),
.B(n_275),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_634),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_735),
.B(n_247),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_815),
.A2(n_803),
.B(n_765),
.C(n_865),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_803),
.A2(n_674),
.B1(n_708),
.B2(n_650),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_772),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_765),
.B(n_650),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_839),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_777),
.B(n_708),
.Y(n_936)
);

CKINVDCx11_ASAP7_75t_R g937 ( 
.A(n_798),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_770),
.B(n_751),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_883),
.A2(n_686),
.B(n_707),
.C(n_753),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_786),
.B(n_704),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_855),
.A2(n_747),
.B1(n_642),
.B2(n_686),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_782),
.B(n_849),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_800),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_830),
.A2(n_756),
.B1(n_763),
.B2(n_714),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_897),
.B(n_656),
.Y(n_945)
);

NOR2x1_ASAP7_75t_L g946 ( 
.A(n_853),
.B(n_653),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_883),
.B(n_451),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_772),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_769),
.A2(n_451),
.B(n_75),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_807),
.A2(n_256),
.B(n_261),
.C(n_263),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_853),
.B(n_841),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_451),
.B(n_70),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_778),
.A2(n_779),
.B(n_790),
.Y(n_953)
);

BUFx4f_ASAP7_75t_L g954 ( 
.A(n_841),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_811),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_790),
.A2(n_65),
.B(n_59),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_841),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_824),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_881),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_831),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_SL g961 ( 
.A1(n_808),
.A2(n_301),
.B1(n_298),
.B2(n_294),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_837),
.B(n_282),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_837),
.B(n_278),
.Y(n_963)
);

BUFx4f_ASAP7_75t_L g964 ( 
.A(n_841),
.Y(n_964)
);

AO21x1_ASAP7_75t_L g965 ( 
.A1(n_920),
.A2(n_247),
.B(n_8),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_837),
.B(n_265),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_781),
.B(n_271),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_812),
.B(n_301),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_781),
.B(n_269),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_847),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_927),
.A2(n_116),
.B(n_77),
.C(n_79),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_930),
.A2(n_140),
.B(n_96),
.C(n_102),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_863),
.B(n_900),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_885),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_863),
.B(n_157),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_878),
.B(n_298),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_804),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_814),
.B(n_294),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_856),
.B(n_290),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_852),
.B(n_290),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_863),
.B(n_147),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_870),
.B(n_286),
.C(n_8),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_825),
.A2(n_7),
.B(n_10),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_790),
.A2(n_144),
.B(n_118),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_790),
.A2(n_108),
.B(n_105),
.Y(n_985)
);

CKINVDCx10_ASAP7_75t_R g986 ( 
.A(n_799),
.Y(n_986)
);

OAI22x1_ASAP7_75t_L g987 ( 
.A1(n_914),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_766),
.A2(n_797),
.B(n_809),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_887),
.B(n_11),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_863),
.Y(n_990)
);

CKINVDCx16_ASAP7_75t_R g991 ( 
.A(n_867),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_851),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_837),
.B(n_74),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_845),
.B(n_104),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_881),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_850),
.B(n_925),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_842),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_784),
.A2(n_14),
.B1(n_15),
.B2(n_21),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_845),
.B(n_881),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_795),
.A2(n_22),
.B(n_23),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_804),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_845),
.B(n_22),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_845),
.B(n_23),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_871),
.B(n_25),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_L g1005 ( 
.A(n_870),
.B(n_25),
.C(n_26),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_917),
.B(n_26),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_919),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_881),
.B(n_27),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_822),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_810),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_838),
.A2(n_44),
.B(n_45),
.Y(n_1011)
);

INVx6_ASAP7_75t_L g1012 ( 
.A(n_821),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_823),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_850),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_794),
.B(n_45),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_825),
.B(n_46),
.Y(n_1016)
);

OA21x2_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_46),
.B(n_48),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_889),
.B(n_52),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_783),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_889),
.B(n_53),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_835),
.B(n_53),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_821),
.A2(n_58),
.B1(n_906),
.B2(n_894),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_867),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_861),
.B(n_846),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_785),
.A2(n_789),
.B(n_788),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_801),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_832),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_909),
.B(n_890),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_854),
.A2(n_771),
.B(n_780),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_774),
.B(n_768),
.Y(n_1030)
);

INVx3_ASAP7_75t_SL g1031 ( 
.A(n_860),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_890),
.B(n_916),
.C(n_872),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_801),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_818),
.B(n_922),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_893),
.B(n_895),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_817),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_773),
.A2(n_872),
.B(n_818),
.C(n_911),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_907),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_925),
.A2(n_859),
.B1(n_869),
.B2(n_926),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_875),
.B(n_926),
.C(n_928),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_899),
.B(n_929),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_848),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_791),
.A2(n_880),
.B(n_857),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_929),
.B(n_775),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_829),
.A2(n_826),
.B(n_792),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_775),
.B(n_857),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_891),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_882),
.B(n_913),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_793),
.B(n_902),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_886),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_891),
.B(n_901),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_886),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_898),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_882),
.B(n_913),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_904),
.B(n_918),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_SL g1056 ( 
.A(n_787),
.B(n_903),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_SL g1057 ( 
.A1(n_816),
.A2(n_833),
.B(n_873),
.C(n_862),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_908),
.B(n_912),
.Y(n_1058)
);

OA22x2_ASAP7_75t_L g1059 ( 
.A1(n_864),
.A2(n_836),
.B1(n_827),
.B2(n_819),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_896),
.B(n_924),
.Y(n_1060)
);

BUFx5_ASAP7_75t_L g1061 ( 
.A(n_813),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_921),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_879),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_843),
.B(n_844),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_840),
.B(n_877),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_820),
.B(n_828),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_874),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_858),
.B(n_888),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_SL g1069 ( 
.A1(n_876),
.A2(n_868),
.B(n_866),
.C(n_884),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_892),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_L g1071 ( 
.A1(n_1016),
.A2(n_910),
.B(n_802),
.C(n_805),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_1018),
.B(n_905),
.C(n_923),
.Y(n_1072)
);

BUFx4_ASAP7_75t_SL g1073 ( 
.A(n_1036),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_953),
.A2(n_796),
.B(n_806),
.Y(n_1074)
);

INVx6_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_988),
.A2(n_915),
.B(n_1025),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_986),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_1050),
.A2(n_1037),
.A3(n_1066),
.B(n_1052),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1065),
.A2(n_1064),
.B(n_1051),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_1030),
.A2(n_965),
.A3(n_1049),
.B(n_1043),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_959),
.B(n_954),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_974),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_SL g1083 ( 
.A1(n_932),
.A2(n_936),
.B(n_1024),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_SL g1084 ( 
.A1(n_998),
.A2(n_983),
.B1(n_1010),
.B2(n_1020),
.C(n_932),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_1045),
.A2(n_1030),
.B(n_952),
.C(n_949),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_955),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_958),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1038),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_1039),
.A2(n_1005),
.B1(n_982),
.B2(n_967),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_960),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_959),
.B(n_954),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_1067),
.A2(n_1024),
.A3(n_1058),
.B(n_1055),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1028),
.A2(n_934),
.B1(n_969),
.B2(n_998),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1069),
.A2(n_1029),
.B(n_1045),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1014),
.B(n_1032),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_939),
.A2(n_1021),
.B(n_1006),
.C(n_978),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_968),
.A2(n_978),
.B(n_989),
.C(n_1008),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_950),
.A2(n_1046),
.B(n_1040),
.C(n_936),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_970),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1014),
.B(n_948),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_964),
.Y(n_1101)
);

OAI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_961),
.A2(n_976),
.B1(n_941),
.B2(n_1022),
.C(n_1009),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_977),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_1070),
.A2(n_1053),
.A3(n_947),
.B(n_987),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_992),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1001),
.Y(n_1106)
);

O2A1O1Ixp5_ASAP7_75t_SL g1107 ( 
.A1(n_1002),
.A2(n_1003),
.B(n_962),
.C(n_966),
.Y(n_1107)
);

OAI22x1_ASAP7_75t_L g1108 ( 
.A1(n_948),
.A2(n_1017),
.B1(n_996),
.B2(n_1015),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_996),
.A2(n_1012),
.B1(n_940),
.B2(n_1014),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1056),
.A2(n_1068),
.B(n_942),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1059),
.A2(n_1057),
.B(n_1011),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1013),
.B(n_1027),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1000),
.A2(n_938),
.A3(n_1004),
.B(n_1042),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1019),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_945),
.Y(n_1115)
);

AO21x1_ASAP7_75t_L g1116 ( 
.A1(n_1068),
.A2(n_1048),
.B(n_1054),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_968),
.A2(n_963),
.B(n_979),
.C(n_980),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1041),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1047),
.A2(n_1035),
.B(n_946),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_979),
.A2(n_980),
.B(n_1007),
.C(n_994),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1060),
.A2(n_945),
.B(n_999),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1023),
.B(n_1012),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1063),
.A2(n_1044),
.B(n_959),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_973),
.B(n_997),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_971),
.A2(n_972),
.B(n_944),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1063),
.A2(n_959),
.B(n_1033),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_964),
.B(n_951),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_951),
.B(n_990),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_956),
.A2(n_985),
.A3(n_984),
.B(n_1017),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_937),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_993),
.A2(n_995),
.B(n_981),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_993),
.B(n_975),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1062),
.A2(n_975),
.B1(n_981),
.B2(n_1019),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1031),
.A2(n_935),
.B(n_1062),
.C(n_1061),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1026),
.A2(n_990),
.A3(n_1061),
.B(n_1019),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_957),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_957),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1061),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1028),
.B(n_624),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_932),
.A2(n_803),
.B1(n_647),
.B2(n_784),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_957),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_931),
.A2(n_803),
.B(n_815),
.C(n_647),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_931),
.A2(n_803),
.B(n_815),
.C(n_647),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1034),
.A2(n_815),
.B(n_1037),
.C(n_865),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_1018),
.A2(n_1020),
.B1(n_1016),
.B2(n_803),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_948),
.B(n_767),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1028),
.B(n_803),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_991),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_974),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_934),
.B(n_803),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_931),
.A2(n_815),
.B(n_803),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_986),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1016),
.A2(n_765),
.B(n_1018),
.Y(n_1153)
);

INVx6_ASAP7_75t_L g1154 ( 
.A(n_991),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1028),
.B(n_803),
.Y(n_1156)
);

OR2x6_ASAP7_75t_SL g1157 ( 
.A(n_1023),
.B(n_506),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_803),
.Y(n_1158)
);

AOI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1018),
.A2(n_765),
.B1(n_666),
.B2(n_1020),
.C(n_1016),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1028),
.B(n_803),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_996),
.B(n_951),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1016),
.A2(n_803),
.B1(n_765),
.B2(n_1018),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1028),
.B(n_624),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1016),
.A2(n_815),
.B(n_647),
.C(n_803),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_1041),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1167)
);

OA22x2_ASAP7_75t_L g1168 ( 
.A1(n_987),
.A2(n_396),
.B1(n_480),
.B2(n_470),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_986),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_986),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_815),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_934),
.B(n_803),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_931),
.A2(n_815),
.B(n_803),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_943),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_1050),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_954),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_954),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_933),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_L g1181 ( 
.A(n_1032),
.B(n_815),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_815),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_953),
.A2(n_554),
.B(n_525),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_1050),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1025),
.A2(n_815),
.A3(n_1050),
.B(n_768),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1028),
.B(n_803),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_931),
.A2(n_803),
.B(n_815),
.C(n_647),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1028),
.B(n_647),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_943),
.Y(n_1191)
);

AND2x6_ASAP7_75t_SL g1192 ( 
.A(n_1016),
.B(n_1018),
.Y(n_1192)
);

AOI221x1_ASAP7_75t_L g1193 ( 
.A1(n_1016),
.A2(n_815),
.B1(n_803),
.B2(n_1020),
.C(n_1018),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1028),
.B(n_803),
.Y(n_1194)
);

OAI22x1_ASAP7_75t_L g1195 ( 
.A1(n_1018),
.A2(n_1020),
.B1(n_1016),
.B2(n_803),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_931),
.A2(n_815),
.B(n_803),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1140),
.A2(n_1168),
.B1(n_1102),
.B2(n_1181),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1146),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1077),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1087),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1150),
.B(n_1173),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1176),
.Y(n_1202)
);

BUFx2_ASAP7_75t_SL g1203 ( 
.A(n_1172),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_1162),
.B2(n_1145),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1153),
.A2(n_1162),
.B1(n_1195),
.B2(n_1089),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1093),
.A2(n_1140),
.B1(n_1151),
.B2(n_1196),
.Y(n_1206)
);

BUFx2_ASAP7_75t_SL g1207 ( 
.A(n_1172),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1086),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1151),
.A2(n_1196),
.B1(n_1174),
.B2(n_1190),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1093),
.A2(n_1143),
.B1(n_1189),
.B2(n_1142),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1174),
.A2(n_1184),
.B1(n_1171),
.B2(n_1192),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1193),
.A2(n_1147),
.B1(n_1188),
.B2(n_1194),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1150),
.B(n_1173),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1172),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1090),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1179),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1141),
.B(n_1178),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1130),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1178),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1112),
.A2(n_1164),
.B1(n_1158),
.B2(n_1156),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1099),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1105),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1096),
.A2(n_1097),
.B(n_1118),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1117),
.A2(n_1163),
.B(n_1139),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1157),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1171),
.A2(n_1184),
.B1(n_1160),
.B2(n_1095),
.Y(n_1226)
);

BUFx8_ASAP7_75t_SL g1227 ( 
.A(n_1152),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_1179),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1169),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1149),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1081),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1116),
.A2(n_1132),
.B1(n_1110),
.B2(n_1192),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1084),
.A2(n_1154),
.B1(n_1075),
.B2(n_1112),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1133),
.A2(n_1115),
.B1(n_1083),
.B2(n_1191),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1109),
.A2(n_1098),
.B(n_1120),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1075),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1141),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

BUFx4f_ASAP7_75t_SL g1239 ( 
.A(n_1148),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1154),
.A2(n_1124),
.B1(n_1161),
.B2(n_1088),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1081),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1103),
.Y(n_1242)
);

INVx6_ASAP7_75t_L g1243 ( 
.A(n_1128),
.Y(n_1243)
);

BUFx8_ASAP7_75t_L g1244 ( 
.A(n_1082),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1100),
.A2(n_1165),
.B1(n_1108),
.B2(n_1115),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1170),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1078),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1084),
.A2(n_1122),
.B1(n_1165),
.B2(n_1144),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1078),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1180),
.A2(n_1131),
.B1(n_1101),
.B2(n_1121),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_SL g1251 ( 
.A(n_1137),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1079),
.A2(n_1177),
.B1(n_1186),
.B2(n_1091),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1114),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1072),
.A2(n_1125),
.B1(n_1138),
.B2(n_1123),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1094),
.A2(n_1127),
.B1(n_1111),
.B2(n_1091),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1113),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1073),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1134),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1076),
.A2(n_1136),
.B1(n_1119),
.B2(n_1126),
.Y(n_1259)
);

INVx3_ASAP7_75t_SL g1260 ( 
.A(n_1107),
.Y(n_1260)
);

BUFx10_ASAP7_75t_L g1261 ( 
.A(n_1135),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1085),
.A2(n_1155),
.B1(n_1185),
.B2(n_1167),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1104),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1166),
.A2(n_1182),
.B1(n_1175),
.B2(n_1183),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1074),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1104),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1080),
.Y(n_1267)
);

OAI22x1_ASAP7_75t_L g1268 ( 
.A1(n_1092),
.A2(n_1080),
.B1(n_1187),
.B2(n_1129),
.Y(n_1268)
);

BUFx4f_ASAP7_75t_SL g1269 ( 
.A(n_1187),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1080),
.B(n_1129),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1129),
.A2(n_998),
.B1(n_803),
.B2(n_932),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1071),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1140),
.A2(n_998),
.B1(n_803),
.B2(n_932),
.Y(n_1273)
);

CKINVDCx11_ASAP7_75t_R g1274 ( 
.A(n_1157),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1162),
.A2(n_647),
.B1(n_1193),
.B2(n_1159),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1146),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1172),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1193),
.A2(n_815),
.B(n_803),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_1162),
.B2(n_803),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1087),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1162),
.A2(n_932),
.B1(n_1159),
.B2(n_1153),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1162),
.A2(n_647),
.B1(n_1193),
.B2(n_1159),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1161),
.B(n_1178),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1073),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1087),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1087),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1141),
.B(n_1178),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1162),
.A2(n_647),
.B1(n_1193),
.B2(n_1159),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1162),
.A2(n_647),
.B1(n_1193),
.B2(n_1159),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1087),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1178),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1157),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_803),
.B2(n_1162),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1077),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_803),
.B2(n_1162),
.Y(n_1296)
);

CKINVDCx6p67_ASAP7_75t_R g1297 ( 
.A(n_1149),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1087),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_1148),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1192),
.B(n_1153),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1140),
.A2(n_998),
.B1(n_803),
.B2(n_932),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_1162),
.B2(n_803),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1172),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_803),
.B2(n_1162),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1148),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1162),
.A2(n_932),
.B1(n_1159),
.B2(n_1153),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1157),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_803),
.B2(n_1162),
.Y(n_1308)
);

INVx6_ASAP7_75t_L g1309 ( 
.A(n_1178),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1148),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1150),
.B(n_1173),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1210),
.B(n_1264),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1256),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1210),
.B(n_1272),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1247),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1211),
.B(n_1209),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1249),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1227),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1199),
.Y(n_1320)
);

OAI21xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1206),
.A2(n_1302),
.B(n_1279),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1201),
.B(n_1213),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1267),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1201),
.B(n_1213),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1211),
.B(n_1209),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1305),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1270),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1268),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1198),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1269),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1261),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1311),
.B(n_1276),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1208),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1265),
.B(n_1259),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1215),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1221),
.Y(n_1336)
);

INVx8_ASAP7_75t_L g1337 ( 
.A(n_1251),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1226),
.B(n_1197),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1222),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1311),
.B(n_1220),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1238),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1263),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1252),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1197),
.B(n_1205),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1278),
.B(n_1271),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1252),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1254),
.A2(n_1235),
.B(n_1223),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1220),
.A2(n_1281),
.B(n_1306),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1271),
.B(n_1204),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1250),
.B(n_1231),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1242),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1273),
.B(n_1301),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1200),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1202),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1231),
.B(n_1280),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1253),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1285),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1286),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1291),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1273),
.B(n_1301),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1298),
.Y(n_1361)
);

AO21x1_ASAP7_75t_L g1362 ( 
.A1(n_1275),
.A2(n_1289),
.B(n_1288),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1281),
.A2(n_1306),
.B(n_1234),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1234),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1255),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1260),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_SL g1367 ( 
.A(n_1219),
.B(n_1292),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1260),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1255),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1262),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1262),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1275),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1282),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1258),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1282),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1241),
.B(n_1248),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1232),
.A2(n_1245),
.B(n_1308),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1212),
.B(n_1296),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1294),
.A2(n_1304),
.B(n_1224),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1217),
.A2(n_1287),
.B(n_1240),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1300),
.A2(n_1289),
.B(n_1288),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1233),
.A2(n_1309),
.B1(n_1292),
.B2(n_1219),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1292),
.B(n_1309),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1233),
.A2(n_1309),
.B1(n_1236),
.B2(n_1243),
.Y(n_1384)
);

INVx5_ASAP7_75t_L g1385 ( 
.A(n_1243),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1217),
.A2(n_1237),
.B(n_1243),
.Y(n_1386)
);

AOI211xp5_ASAP7_75t_L g1387 ( 
.A1(n_1257),
.A2(n_1230),
.B(n_1284),
.C(n_1283),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_1299),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1277),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1388),
.B(n_1239),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1388),
.B(n_1310),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1321),
.A2(n_1228),
.B(n_1216),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1321),
.A2(n_1307),
.B1(n_1274),
.B2(n_1293),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1379),
.A2(n_1203),
.B(n_1207),
.C(n_1303),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1322),
.B(n_1214),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1329),
.B(n_1297),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1379),
.A2(n_1225),
.B(n_1277),
.C(n_1251),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1330),
.B(n_1228),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_SL g1399 ( 
.A1(n_1387),
.A2(n_1244),
.B(n_1229),
.C(n_1199),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1363),
.A2(n_1244),
.B(n_1246),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1342),
.B(n_1246),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1342),
.B(n_1295),
.Y(n_1402)
);

AND2x6_ASAP7_75t_L g1403 ( 
.A(n_1352),
.B(n_1218),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1362),
.A2(n_1290),
.B1(n_1295),
.B2(n_1344),
.Y(n_1404)
);

NAND2x1_ASAP7_75t_L g1405 ( 
.A(n_1367),
.B(n_1383),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1351),
.B(n_1341),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1319),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1362),
.A2(n_1352),
.B1(n_1360),
.B2(n_1344),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1330),
.B(n_1350),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1333),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1324),
.B(n_1332),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1360),
.A2(n_1377),
.B(n_1349),
.C(n_1378),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1333),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1364),
.A2(n_1384),
.B(n_1312),
.C(n_1349),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1377),
.A2(n_1345),
.B(n_1338),
.C(n_1325),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1350),
.B(n_1355),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1326),
.B(n_1374),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1312),
.A2(n_1340),
.B(n_1375),
.C(n_1373),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1317),
.A2(n_1325),
.B(n_1334),
.C(n_1375),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1335),
.B(n_1339),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1334),
.A2(n_1372),
.B(n_1371),
.C(n_1370),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1356),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1343),
.A2(n_1346),
.B(n_1368),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1348),
.A2(n_1347),
.B(n_1381),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1353),
.B(n_1354),
.Y(n_1426)
);

NAND2x1_ASAP7_75t_L g1427 ( 
.A(n_1367),
.B(n_1383),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1337),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_R g1429 ( 
.A(n_1347),
.B(n_1381),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1355),
.B(n_1334),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1355),
.B(n_1350),
.Y(n_1431)
);

AO32x1_ASAP7_75t_L g1432 ( 
.A1(n_1366),
.A2(n_1368),
.A3(n_1328),
.B1(n_1382),
.B2(n_1323),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_SL g1433 ( 
.A(n_1312),
.B(n_1314),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1380),
.A2(n_1387),
.B(n_1337),
.C(n_1369),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1374),
.B(n_1320),
.Y(n_1435)
);

NAND4xp25_ASAP7_75t_L g1436 ( 
.A(n_1358),
.B(n_1359),
.C(n_1361),
.D(n_1366),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1353),
.B(n_1354),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1357),
.B(n_1336),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1380),
.A2(n_1337),
.B(n_1365),
.C(n_1369),
.Y(n_1439)
);

OAI211xp5_ASAP7_75t_L g1440 ( 
.A1(n_1365),
.A2(n_1328),
.B(n_1374),
.C(n_1346),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1314),
.A2(n_1376),
.B(n_1386),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1424),
.B(n_1327),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1424),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1410),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1413),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1421),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1425),
.B(n_1313),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1437),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1418),
.A2(n_1374),
.B1(n_1337),
.B2(n_1385),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1438),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1406),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1431),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1416),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1409),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1436),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1433),
.B(n_1315),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1441),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1436),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1405),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1423),
.B(n_1316),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1461),
.B(n_1458),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1454),
.B(n_1430),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1446),
.A2(n_1404),
.B1(n_1408),
.B2(n_1393),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1446),
.A2(n_1393),
.B1(n_1429),
.B2(n_1412),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1443),
.B(n_1440),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1423),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1459),
.B(n_1427),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1444),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1457),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1415),
.Y(n_1473)
);

AOI221x1_ASAP7_75t_L g1474 ( 
.A1(n_1457),
.A2(n_1394),
.B1(n_1397),
.B2(n_1420),
.C(n_1400),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1454),
.B(n_1439),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1454),
.B(n_1316),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1457),
.A2(n_1434),
.B1(n_1414),
.B2(n_1422),
.C(n_1400),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1460),
.A2(n_1419),
.B1(n_1392),
.B2(n_1395),
.C(n_1411),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1453),
.B(n_1390),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1460),
.A2(n_1399),
.B1(n_1391),
.B2(n_1435),
.C(n_1417),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1453),
.B(n_1401),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1455),
.B(n_1402),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1445),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1445),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1452),
.B(n_1318),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1448),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1445),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1455),
.B(n_1331),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1461),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1463),
.B(n_1461),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1475),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1484),
.Y(n_1495)
);

NAND3x1_ASAP7_75t_SL g1496 ( 
.A(n_1474),
.B(n_1403),
.C(n_1432),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1484),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1473),
.B(n_1453),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1485),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1463),
.B(n_1459),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1475),
.B(n_1459),
.Y(n_1501)
);

CKINVDCx16_ASAP7_75t_R g1502 ( 
.A(n_1467),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1471),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1455),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1468),
.B(n_1473),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1485),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1469),
.B(n_1460),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1487),
.B(n_1462),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1470),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1489),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1489),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1477),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1477),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1477),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1470),
.B(n_1461),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1470),
.B(n_1461),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1503),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1502),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1506),
.B(n_1479),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1495),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1503),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1495),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1497),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1535)
);

AND2x4_ASAP7_75t_SL g1536 ( 
.A(n_1491),
.B(n_1428),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1499),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1498),
.B(n_1479),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1509),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1498),
.B(n_1469),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1483),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1505),
.B(n_1511),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1483),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1514),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1513),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1514),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1505),
.B(n_1465),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1465),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1492),
.B(n_1476),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1491),
.B(n_1490),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_SL g1556 ( 
.A(n_1513),
.B(n_1456),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1492),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1501),
.B(n_1476),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1508),
.B(n_1521),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.B(n_1521),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1526),
.Y(n_1562)
);

AND2x2_ASAP7_75t_SL g1563 ( 
.A(n_1524),
.B(n_1466),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1551),
.B(n_1516),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1524),
.B(n_1481),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1551),
.B(n_1517),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1541),
.B(n_1517),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1556),
.B(n_1513),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1541),
.B(n_1550),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1535),
.B(n_1493),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1535),
.B(n_1493),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1480),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1493),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1545),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1526),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1493),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1529),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1482),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1529),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1530),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1530),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1519),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1525),
.A2(n_1467),
.B(n_1466),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1523),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1539),
.B(n_1504),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1539),
.B(n_1544),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1550),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1523),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1531),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1544),
.B(n_1481),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1536),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1534),
.B(n_1519),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1561),
.B(n_1512),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1534),
.B(n_1519),
.Y(n_1597)
);

NAND2x1p5_ASAP7_75t_L g1598 ( 
.A(n_1591),
.B(n_1563),
.Y(n_1598)
);

OAI321xp33_ASAP7_75t_L g1599 ( 
.A1(n_1584),
.A2(n_1548),
.A3(n_1478),
.B1(n_1534),
.B2(n_1522),
.C(n_1558),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1565),
.A2(n_1548),
.B(n_1478),
.C(n_1558),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1562),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1563),
.A2(n_1556),
.B(n_1474),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1570),
.Y(n_1605)
);

AOI21xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1563),
.A2(n_1548),
.B(n_1407),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1568),
.Y(n_1607)
);

NAND3x2_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1522),
.C(n_1561),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1587),
.A2(n_1396),
.B(n_1554),
.C(n_1557),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1572),
.Y(n_1610)
);

NOR3xp33_ASAP7_75t_SL g1611 ( 
.A(n_1578),
.B(n_1554),
.C(n_1537),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1568),
.A2(n_1528),
.B(n_1523),
.Y(n_1612)
);

XNOR2xp5_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1389),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1593),
.A2(n_1597),
.B1(n_1574),
.B2(n_1586),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1574),
.B(n_1536),
.Y(n_1616)
);

OAI32xp33_ASAP7_75t_L g1617 ( 
.A1(n_1588),
.A2(n_1496),
.A3(n_1532),
.B1(n_1527),
.B2(n_1559),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1575),
.Y(n_1618)
);

OAI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1583),
.A2(n_1569),
.B1(n_1513),
.B2(n_1566),
.C(n_1564),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1569),
.Y(n_1620)
);

AOI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1564),
.A2(n_1513),
.B(n_1531),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1577),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1571),
.B(n_1555),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1601),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1612),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1598),
.A2(n_1579),
.B(n_1577),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1598),
.A2(n_1580),
.B(n_1579),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1603),
.B(n_1580),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1598),
.A2(n_1616),
.B1(n_1608),
.B2(n_1615),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1599),
.B(n_1513),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1604),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1597),
.B1(n_1593),
.B2(n_1582),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1611),
.B(n_1590),
.C(n_1581),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1607),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1618),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1622),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1581),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1613),
.B(n_1582),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1605),
.Y(n_1642)
);

AOI221x1_ASAP7_75t_L g1643 ( 
.A1(n_1626),
.A2(n_1606),
.B1(n_1621),
.B2(n_1615),
.C(n_1605),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1628),
.B(n_1600),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1637),
.B(n_1614),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1625),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1637),
.Y(n_1647)
);

NAND3x2_ASAP7_75t_L g1648 ( 
.A(n_1642),
.B(n_1608),
.C(n_1624),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1641),
.B(n_1573),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1631),
.A2(n_1613),
.B1(n_1619),
.B2(n_1623),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_L g1651 ( 
.A1(n_1629),
.A2(n_1617),
.B(n_1573),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1633),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1636),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_L g1654 ( 
.A(n_1652),
.B(n_1640),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1644),
.B(n_1640),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1634),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1643),
.B(n_1626),
.C(n_1627),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1658)
);

NAND2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1647),
.B(n_1630),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1648),
.B(n_1638),
.C(n_1632),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1653),
.B(n_1639),
.C(n_1609),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1651),
.A2(n_1590),
.B(n_1566),
.C(n_1576),
.Y(n_1663)
);

NOR3x1_ASAP7_75t_L g1664 ( 
.A(n_1657),
.B(n_1650),
.C(n_1645),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1655),
.A2(n_1649),
.B1(n_1646),
.B2(n_1536),
.Y(n_1665)
);

OAI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1658),
.A2(n_1646),
.B(n_1649),
.C(n_1612),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1656),
.A2(n_1576),
.B1(n_1585),
.B2(n_1589),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1659),
.Y(n_1668)
);

AOI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1660),
.A2(n_1612),
.B(n_1589),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1661),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_SL g1671 ( 
.A(n_1668),
.B(n_1663),
.C(n_1662),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1666),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1670),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1654),
.B(n_1389),
.C(n_1585),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1667),
.A2(n_1596),
.B1(n_1567),
.B2(n_1594),
.C(n_1595),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1669),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1664),
.A2(n_1596),
.B1(n_1567),
.B2(n_1594),
.C(n_1595),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1673),
.Y(n_1678)
);

AOI31xp33_ASAP7_75t_L g1679 ( 
.A1(n_1674),
.A2(n_1451),
.A3(n_1519),
.B(n_1520),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1676),
.Y(n_1680)
);

NOR2x1_ASAP7_75t_L g1681 ( 
.A(n_1671),
.B(n_1537),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1538),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1678),
.A2(n_1681),
.B(n_1679),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_L g1684 ( 
.A(n_1680),
.B(n_1677),
.C(n_1675),
.Y(n_1684)
);

OAI321xp33_ASAP7_75t_L g1685 ( 
.A1(n_1682),
.A2(n_1532),
.A3(n_1527),
.B1(n_1533),
.B2(n_1528),
.C(n_1553),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1684),
.B(n_1451),
.C(n_1428),
.D(n_1520),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1686),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1687),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1687),
.A2(n_1683),
.B(n_1685),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1689),
.A2(n_1528),
.B1(n_1533),
.B2(n_1553),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1690),
.A2(n_1688),
.B1(n_1533),
.B2(n_1540),
.Y(n_1692)
);

AO21x1_ASAP7_75t_L g1693 ( 
.A1(n_1691),
.A2(n_1553),
.B(n_1540),
.Y(n_1693)
);

CKINVDCx16_ASAP7_75t_R g1694 ( 
.A(n_1692),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1693),
.B(n_1540),
.Y(n_1695)
);

XOR2xp5_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1398),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1552),
.B1(n_1538),
.B2(n_1557),
.C(n_1542),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1549),
.B(n_1546),
.C(n_1547),
.Y(n_1698)
);


endmodule