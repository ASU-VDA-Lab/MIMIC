module fake_aes_9581_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
AND2x6_ASAP7_75t_L g15 ( .A(n_8), .B(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_2), .Y(n_19) );
BUFx5_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_16), .B(n_13), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_17), .Y(n_23) );
OAI21x1_ASAP7_75t_L g24 ( .A1(n_19), .A2(n_12), .B(n_15), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_22), .Y(n_26) );
INVx2_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_25), .B(n_23), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_28), .B(n_23), .Y(n_29) );
OAI32xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_26), .A3(n_15), .B1(n_24), .B2(n_2), .Y(n_30) );
AOI21xp33_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_3), .B(n_4), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OAI221xp5_ASAP7_75t_SL g33 ( .A1(n_30), .A2(n_26), .B1(n_15), .B2(n_3), .C(n_24), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_32), .B(n_15), .Y(n_34) );
NAND2xp33_ASAP7_75t_SL g35 ( .A(n_32), .B(n_5), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_31), .Y(n_36) );
NOR4xp25_ASAP7_75t_L g37 ( .A(n_36), .B(n_33), .C(n_9), .D(n_10), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
OR2x2_ASAP7_75t_L g39 ( .A(n_38), .B(n_35), .Y(n_39) );
OA22x2_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_37), .B1(n_7), .B2(n_20), .Y(n_40) );
endmodule