module real_jpeg_5366_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_3),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_3),
.B(n_207),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_4),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_4),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_4),
.B(n_35),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_4),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_4),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_5),
.B(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_7),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_8),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_8),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_35),
.Y(n_242)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_10),
.Y(n_176)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_11),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_13),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_13),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_13),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_30),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

AND2x6_ASAP7_75t_SL g183 ( 
.A(n_16),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_16),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_16),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_16),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_16),
.B(n_52),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_16),
.B(n_276),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_17),
.Y(n_154)
);

XNOR2x2_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_194),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_193),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_164),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_22),
.B(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_93),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_62),
.C(n_75),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_24),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.C(n_49),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_25),
.A2(n_26),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_27),
.B(n_33),
.C(n_40),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_28),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_42),
.B(n_50),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_43),
.B(n_46),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_45),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_45),
.Y(n_173)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_45),
.Y(n_205)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_48),
.Y(n_216)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_60),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_51),
.B(n_60),
.Y(n_289)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_55),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_57),
.Y(n_249)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_58),
.Y(n_273)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_59),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_61),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_62),
.B(n_75),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_68),
.C(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_86),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_82),
.C(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_81),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_81),
.Y(n_254)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_86),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.C(n_90),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_89),
.Y(n_189)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_125),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_146),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_145),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_127),
.A2(n_128),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_132),
.C(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_162),
.B2(n_163),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_190),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_166),
.B(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_168),
.B(n_190),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_185),
.C(n_186),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_169),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.C(n_182),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_170),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_266)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_SL g285 ( 
.A(n_178),
.B(n_183),
.Y(n_285)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

AOI21x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_310),
.B(n_314),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_297),
.B(n_309),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_281),
.B(n_296),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_257),
.B(n_280),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_238),
.B(n_256),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_218),
.B(n_237),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_212),
.B(n_217),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_209),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_206),
.Y(n_219)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_229),
.C(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_255),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_255),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_244),
.C(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_269),
.C(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_260),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_268),
.C(n_271),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_277),
.C(n_278),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_295),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_286),
.C(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_292),
.C(n_293),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_307),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.C(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_313),
.Y(n_314)
);


endmodule