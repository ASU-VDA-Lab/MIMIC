module fake_ariane_2934_n_1117 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1117);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1117;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_1018;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_770;
wire n_928;
wire n_839;
wire n_1099;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_847;
wire n_747;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_998;
wire n_999;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_1069;
wire n_965;
wire n_393;
wire n_886;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_117),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_171),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_1),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_84),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_91),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_65),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_103),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_69),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_85),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_167),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_61),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_51),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_72),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_123),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_199),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_147),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_66),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_73),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_55),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_46),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_14),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_160),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_188),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_93),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_78),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_185),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_150),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_74),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_10),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_166),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_172),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_226),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_263),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_231),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_217),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_223),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_220),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_207),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_207),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_257),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_234),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_234),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_253),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_258),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_258),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_261),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_291),
.A2(n_257),
.B(n_210),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_216),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_R g331 ( 
.A1(n_316),
.A2(n_324),
.B1(n_325),
.B2(n_323),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_277),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_208),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_211),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_218),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_219),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_227),
.B(n_222),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_316),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_213),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_228),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_230),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_307),
.A2(n_319),
.B1(n_312),
.B2(n_285),
.Y(n_354)
);

CKINVDCx6p67_ASAP7_75t_R g355 ( 
.A(n_285),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_232),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_281),
.B(n_213),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_213),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_262),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_236),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_300),
.B(n_237),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_262),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_324),
.B(n_241),
.Y(n_381)
);

AOI22x1_ASAP7_75t_SL g382 ( 
.A1(n_312),
.A2(n_278),
.B1(n_275),
.B2(n_272),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

AO22x2_ASAP7_75t_L g386 ( 
.A1(n_370),
.A2(n_319),
.B1(n_322),
.B2(n_325),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_244),
.C(n_243),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_332),
.B(n_326),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_340),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_246),
.Y(n_404)
);

AND3x2_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_326),
.C(n_0),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_247),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_347),
.B(n_248),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_249),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_250),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_361),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_367),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_256),
.Y(n_418)
);

NOR2x1p5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_260),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

AND3x2_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_1),
.C(n_2),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_332),
.A2(n_271),
.B1(n_270),
.B2(n_267),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_L g428 ( 
.A(n_380),
.B(n_374),
.Y(n_428)
);

OA22x2_ASAP7_75t_L g429 ( 
.A1(n_360),
.A2(n_266),
.B1(n_3),
.B2(n_4),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_359),
.Y(n_433)
);

NOR2x1p5_ASAP7_75t_L g434 ( 
.A(n_380),
.B(n_2),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_329),
.A2(n_35),
.B(n_34),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_36),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_365),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_332),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_345),
.B(n_5),
.C(n_6),
.Y(n_449)
);

BUFx6f_ASAP7_75t_SL g450 ( 
.A(n_377),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_346),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_348),
.Y(n_454)
);

AO21x2_ASAP7_75t_L g455 ( 
.A1(n_358),
.A2(n_38),
.B(n_37),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_6),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_374),
.B(n_7),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_329),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_378),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_378),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_395),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_432),
.B(n_380),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_442),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_454),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_379),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_392),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_420),
.B(n_347),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_372),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_450),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_432),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_412),
.B(n_374),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_420),
.B(n_347),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_375),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_386),
.B(n_370),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_386),
.B(n_348),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_450),
.B(n_405),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_386),
.B(n_354),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_432),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_442),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_432),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_443),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_385),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_386),
.B(n_382),
.Y(n_508)
);

BUFx8_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_443),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_441),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_385),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_448),
.B(n_376),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_406),
.B(n_330),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_SL g519 ( 
.A(n_419),
.B(n_374),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_416),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_446),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_419),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_456),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_456),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_449),
.B(n_377),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_388),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_421),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_423),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_400),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_445),
.B(n_374),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_445),
.B(n_377),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_446),
.B(n_382),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_424),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_430),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_434),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_476),
.A2(n_429),
.B1(n_449),
.B2(n_331),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_409),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_491),
.B(n_451),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_491),
.B(n_451),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_533),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_459),
.B(n_404),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_461),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_462),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_474),
.Y(n_554)
);

O2A1O1Ixp5_ASAP7_75t_L g555 ( 
.A1(n_465),
.A2(n_457),
.B(n_453),
.C(n_437),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_513),
.B(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_513),
.B(n_452),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_460),
.B(n_404),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_460),
.B(n_410),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_355),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_488),
.B(n_476),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_480),
.B(n_355),
.Y(n_563)
);

OAI221xp5_ASAP7_75t_L g564 ( 
.A1(n_498),
.A2(n_373),
.B1(n_356),
.B2(n_410),
.C(n_418),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_468),
.A2(n_452),
.B1(n_429),
.B2(n_418),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_470),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

NAND2x1_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_393),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_497),
.B(n_331),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_504),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_475),
.B(n_400),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_475),
.B(n_400),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_515),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_490),
.B(n_369),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_467),
.B(n_334),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_504),
.B(n_336),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_525),
.A2(n_429),
.B1(n_435),
.B2(n_439),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_517),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_506),
.B(n_435),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_490),
.A2(n_529),
.B1(n_483),
.B2(n_534),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_506),
.B(n_351),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_510),
.B(n_342),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_500),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_510),
.B(n_431),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_519),
.A2(n_428),
.B1(n_434),
.B2(n_350),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_518),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_469),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_536),
.A2(n_431),
.B1(n_439),
.B2(n_433),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_486),
.B(n_433),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_503),
.B(n_400),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_497),
.B(n_371),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_481),
.B(n_356),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_478),
.Y(n_595)
);

NAND2x1_ASAP7_75t_L g596 ( 
.A(n_521),
.B(n_393),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_509),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_499),
.B(n_368),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_369),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_463),
.B(n_369),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_464),
.B(n_390),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_519),
.A2(n_397),
.B1(n_407),
.B2(n_393),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_489),
.B(n_390),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_492),
.B(n_368),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_544),
.B(n_425),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_473),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_493),
.B(n_494),
.Y(n_609)
);

AND2x6_ASAP7_75t_SL g610 ( 
.A(n_495),
.B(n_368),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_505),
.B(n_400),
.Y(n_611)
);

AND2x6_ASAP7_75t_SL g612 ( 
.A(n_508),
.B(n_422),
.Y(n_612)
);

AO22x1_ASAP7_75t_L g613 ( 
.A1(n_509),
.A2(n_458),
.B1(n_438),
.B2(n_453),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_496),
.B(n_425),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_549),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_566),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_554),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_574),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_581),
.B(n_526),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_546),
.B(n_465),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_599),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_549),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_553),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_594),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_579),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_556),
.B(n_477),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_584),
.B(n_553),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_SL g631 ( 
.A(n_593),
.B(n_387),
.C(n_501),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_551),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_567),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_L g635 ( 
.A1(n_587),
.A2(n_502),
.B1(n_345),
.B2(n_533),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_593),
.B(n_524),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_568),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_458),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_569),
.B(n_522),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_550),
.A2(n_425),
.B(n_437),
.C(n_444),
.Y(n_641)
);

AOI21xp33_ASAP7_75t_L g642 ( 
.A1(n_545),
.A2(n_345),
.B(n_531),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_596),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_569),
.A2(n_523),
.B1(n_329),
.B2(n_387),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_561),
.B(n_437),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_SL g646 ( 
.A(n_564),
.B(n_403),
.C(n_402),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_570),
.B(n_583),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_584),
.B(n_417),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_SL g650 ( 
.A(n_588),
.B(n_403),
.C(n_402),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_595),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_608),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_582),
.B(n_543),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_444),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_562),
.B(n_532),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_607),
.Y(n_657)
);

AOI221xp5_ASAP7_75t_SL g658 ( 
.A1(n_545),
.A2(n_444),
.B1(n_541),
.B2(n_540),
.C(n_539),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_558),
.B(n_542),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_590),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_559),
.B(n_537),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_580),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_614),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_585),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_612),
.B(n_397),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_603),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_538),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_605),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_547),
.B(n_484),
.Y(n_671)
);

AOI211xp5_ASAP7_75t_L g672 ( 
.A1(n_565),
.A2(n_414),
.B(n_438),
.C(n_413),
.Y(n_672)
);

AND2x4_ASAP7_75t_SL g673 ( 
.A(n_589),
.B(n_397),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_589),
.B(n_577),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_607),
.B(n_407),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_575),
.B(n_407),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_601),
.B(n_413),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_606),
.Y(n_678)
);

AND3x1_ASAP7_75t_SL g679 ( 
.A(n_610),
.B(n_7),
.C(n_8),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_602),
.B(n_413),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_657),
.B(n_578),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_652),
.Y(n_683)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_624),
.B(n_591),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_640),
.B(n_578),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_671),
.A2(n_436),
.B(n_555),
.Y(n_686)
);

AO31x2_ASAP7_75t_L g687 ( 
.A1(n_671),
.A2(n_557),
.A3(n_507),
.B(n_484),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_636),
.B(n_485),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_629),
.A2(n_573),
.B(n_571),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_620),
.B(n_485),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_627),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_629),
.B(n_571),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_666),
.A2(n_436),
.B(n_573),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_615),
.B(n_630),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_630),
.B(n_507),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_SL g697 ( 
.A1(n_647),
.A2(n_611),
.B(n_591),
.Y(n_697)
);

OAI21x1_ASAP7_75t_SL g698 ( 
.A1(n_647),
.A2(n_604),
.B(n_414),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_623),
.A2(n_611),
.B(n_514),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_666),
.A2(n_656),
.B(n_668),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_672),
.A2(n_613),
.B(n_455),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_667),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_L g703 ( 
.A1(n_674),
.A2(n_455),
.B(n_512),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_620),
.B(n_512),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_681),
.B(n_514),
.Y(n_705)
);

AOI221x1_ASAP7_75t_L g706 ( 
.A1(n_644),
.A2(n_530),
.B1(n_455),
.B2(n_11),
.C(n_12),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_672),
.A2(n_530),
.B(n_417),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_656),
.A2(n_411),
.B(n_417),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_618),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_653),
.A2(n_417),
.B(n_411),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_616),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_616),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_646),
.A2(n_411),
.B(n_417),
.C(n_11),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_653),
.A2(n_417),
.B(n_411),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_617),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_631),
.B(n_8),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_659),
.B(n_411),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_616),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_625),
.Y(n_719)
);

NAND2x1_ASAP7_75t_SL g720 ( 
.A(n_645),
.B(n_411),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_663),
.B(n_9),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_669),
.A2(n_41),
.B(n_40),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_659),
.B(n_9),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_625),
.B(n_43),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_664),
.A2(n_45),
.B(n_44),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_668),
.A2(n_49),
.B(n_47),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_650),
.B(n_12),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_664),
.A2(n_52),
.B(n_50),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_621),
.B(n_13),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_660),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_635),
.A2(n_54),
.B(n_53),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_628),
.B(n_15),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_632),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_641),
.A2(n_57),
.B(n_56),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_677),
.A2(n_127),
.B(n_203),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_634),
.B(n_17),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_673),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_680),
.A2(n_126),
.B(n_201),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_662),
.A2(n_19),
.B(n_20),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_685),
.A2(n_622),
.B1(n_679),
.B2(n_654),
.Y(n_740)
);

AO22x1_ASAP7_75t_L g741 ( 
.A1(n_739),
.A2(n_651),
.B1(n_655),
.B2(n_678),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_702),
.B(n_619),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_708),
.A2(n_649),
.B(n_670),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_701),
.A2(n_644),
.B(n_675),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_731),
.A2(n_675),
.B(n_642),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_697),
.A2(n_707),
.B(n_693),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_SL g747 ( 
.A1(n_713),
.A2(n_642),
.B(n_657),
.C(n_661),
.Y(n_747)
);

BUFx8_ASAP7_75t_SL g748 ( 
.A(n_692),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_695),
.B(n_625),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_739),
.A2(n_658),
.B(n_676),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_682),
.A2(n_658),
.B1(n_676),
.B2(n_639),
.Y(n_751)
);

AOI31xp67_ASAP7_75t_L g752 ( 
.A1(n_693),
.A2(n_648),
.A3(n_638),
.B(n_633),
.Y(n_752)
);

O2A1O1Ixp5_ASAP7_75t_L g753 ( 
.A1(n_722),
.A2(n_639),
.B(n_665),
.C(n_643),
.Y(n_753)
);

BUFx4f_ASAP7_75t_L g754 ( 
.A(n_712),
.Y(n_754)
);

NOR4xp25_ASAP7_75t_L g755 ( 
.A(n_730),
.B(n_20),
.C(n_21),
.D(n_22),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_727),
.A2(n_639),
.B(n_23),
.C(n_24),
.Y(n_756)
);

AOI21xp33_ASAP7_75t_L g757 ( 
.A1(n_717),
.A2(n_665),
.B(n_643),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_706),
.A2(n_639),
.A3(n_665),
.B(n_643),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_683),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_SL g760 ( 
.A1(n_723),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_689),
.A2(n_637),
.B(n_26),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_710),
.A2(n_637),
.B(n_26),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_716),
.A2(n_738),
.B(n_735),
.C(n_732),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_691),
.Y(n_764)
);

BUFx2_ASAP7_75t_R g765 ( 
.A(n_696),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_686),
.A2(n_637),
.B(n_131),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_694),
.A2(n_700),
.B(n_734),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_715),
.B(n_25),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_714),
.A2(n_27),
.B(n_28),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_728),
.A2(n_132),
.B(n_197),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_721),
.B(n_27),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_712),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_709),
.B(n_28),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_733),
.B(n_29),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_699),
.A2(n_29),
.B(n_30),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_712),
.Y(n_776)
);

AOI221x1_ASAP7_75t_L g777 ( 
.A1(n_698),
.A2(n_703),
.B1(n_729),
.B2(n_699),
.C(n_725),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_726),
.A2(n_133),
.B(n_193),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_719),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_736),
.B(n_30),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_711),
.B(n_31),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_684),
.A2(n_31),
.B(n_32),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_688),
.A2(n_135),
.A3(n_192),
.B(n_58),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_719),
.B(n_59),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_720),
.A2(n_32),
.B(n_33),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_737),
.B(n_33),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_705),
.A2(n_60),
.B(n_63),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_SL g790 ( 
.A(n_711),
.B(n_718),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_703),
.A2(n_204),
.B(n_67),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_724),
.A2(n_64),
.B(n_68),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_718),
.B(n_75),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_737),
.A2(n_76),
.B(n_77),
.C(n_79),
.Y(n_794)
);

AO21x2_ASAP7_75t_L g795 ( 
.A1(n_704),
.A2(n_80),
.B(n_82),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_687),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_687),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_687),
.A2(n_191),
.B(n_86),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_701),
.A2(n_189),
.B(n_87),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_701),
.A2(n_187),
.B(n_88),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_SL g801 ( 
.A(n_702),
.B(n_83),
.Y(n_801)
);

AO31x2_ASAP7_75t_L g802 ( 
.A1(n_706),
.A2(n_89),
.A3(n_92),
.B(n_94),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_739),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_683),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_SL g806 ( 
.A1(n_739),
.A2(n_98),
.B(n_99),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_701),
.A2(n_100),
.B(n_102),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_803),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_780),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_740),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_775),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_776),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_764),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_748),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_781),
.B(n_111),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_754),
.Y(n_816)
);

BUFx8_ASAP7_75t_SL g817 ( 
.A(n_776),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_776),
.Y(n_818)
);

INVx6_ASAP7_75t_L g819 ( 
.A(n_779),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_758),
.Y(n_820)
);

BUFx2_ASAP7_75t_SL g821 ( 
.A(n_742),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_786),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_772),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_779),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_786),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_771),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_765),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_749),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_759),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_746),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_783),
.Y(n_831)
);

BUFx12f_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_115),
.Y(n_833)
);

BUFx12f_ASAP7_75t_L g834 ( 
.A(n_774),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_805),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_752),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_768),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_741),
.B(n_184),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_784),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_839)
);

INVx6_ASAP7_75t_L g840 ( 
.A(n_790),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_799),
.A2(n_120),
.B(n_121),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_755),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_842)
);

CKINVDCx11_ASAP7_75t_R g843 ( 
.A(n_797),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_788),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_744),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_751),
.B(n_136),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_796),
.Y(n_847)
);

BUFx4f_ASAP7_75t_L g848 ( 
.A(n_797),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_801),
.B(n_137),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_750),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

INVx6_ASAP7_75t_L g852 ( 
.A(n_797),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_757),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_743),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_758),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_806),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_766),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_756),
.A2(n_145),
.B(n_148),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_760),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_785),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_787),
.B(n_149),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_794),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_785),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_767),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_792),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_847),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_836),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_808),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_822),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_864),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_830),
.B(n_802),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_854),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_862),
.A2(n_795),
.B1(n_761),
.B2(n_745),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_835),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_820),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_813),
.B(n_802),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_857),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_860),
.A2(n_798),
.B(n_800),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_855),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_857),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_831),
.B(n_802),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_822),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_841),
.A2(n_807),
.B(n_804),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_863),
.B(n_777),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_857),
.B(n_763),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_852),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_809),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_809),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_829),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_822),
.B(n_791),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_823),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_825),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_812),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_837),
.B(n_769),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_838),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_858),
.A2(n_762),
.B(n_747),
.Y(n_896)
);

OA21x2_ASAP7_75t_L g897 ( 
.A1(n_838),
.A2(n_753),
.B(n_789),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_848),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_851),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_843),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_846),
.B(n_778),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_825),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_868),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_900),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_895),
.A2(n_858),
.B1(n_842),
.B2(n_811),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_869),
.B(n_846),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_868),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_869),
.B(n_821),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_887),
.B(n_827),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_887),
.B(n_833),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_874),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_866),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_866),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_888),
.B(n_812),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_900),
.B(n_840),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_876),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_867),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_879),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_870),
.Y(n_922)
);

AO21x2_ASAP7_75t_L g923 ( 
.A1(n_895),
.A2(n_842),
.B(n_826),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_891),
.B(n_876),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_892),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_867),
.A2(n_872),
.B(n_883),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_869),
.B(n_849),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_870),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_891),
.B(n_834),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_869),
.B(n_840),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_878),
.A2(n_770),
.B(n_841),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_889),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_892),
.B(n_818),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_921),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_928),
.B(n_827),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_919),
.B(n_871),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_927),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_924),
.B(n_903),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_927),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_918),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_919),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_871),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_926),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_920),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_920),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_929),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_911),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_906),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_910),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_922),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_913),
.B(n_884),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_905),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_929),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_933),
.B(n_903),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_922),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_918),
.B(n_814),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_928),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_917),
.B(n_894),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_938),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_958),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_935),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_935),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_958),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_958),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_949),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_938),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_944),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_944),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_938),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_938),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_917),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_940),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_957),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_952),
.B(n_925),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_942),
.B(n_925),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_964),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_966),
.B(n_948),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_962),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_961),
.B(n_950),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_963),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_961),
.B(n_965),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_968),
.B(n_959),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_969),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_965),
.B(n_950),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_960),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_943),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_977),
.B(n_964),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_979),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_981),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_953),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_987),
.B(n_974),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_980),
.B(n_974),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_977),
.B(n_964),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_993),
.B(n_977),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_SL g996 ( 
.A(n_992),
.B(n_982),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_988),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_991),
.A2(n_936),
.B1(n_890),
.B2(n_978),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_L g999 ( 
.A1(n_991),
.A2(n_890),
.B1(n_940),
.B2(n_908),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_983),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_1000),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_982),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_996),
.B(n_990),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_997),
.B(n_980),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_985),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_995),
.B(n_985),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_1000),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1000),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_995),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_SL g1011 ( 
.A(n_1001),
.B(n_988),
.C(n_994),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1001),
.B(n_986),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_972),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1008),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_1003),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1009),
.B(n_975),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1004),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_1002),
.Y(n_1018)
);

OAI322xp33_ASAP7_75t_L g1019 ( 
.A1(n_1015),
.A2(n_1006),
.A3(n_1005),
.B1(n_1010),
.B2(n_986),
.C1(n_971),
.C2(n_960),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1013),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_930),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1017),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1014),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_1018),
.Y(n_1024)
);

AO22x1_ASAP7_75t_L g1025 ( 
.A1(n_1012),
.A2(n_1016),
.B1(n_1011),
.B2(n_901),
.Y(n_1025)
);

AOI32xp33_ASAP7_75t_L g1026 ( 
.A1(n_1015),
.A2(n_907),
.A3(n_940),
.B1(n_973),
.B2(n_971),
.Y(n_1026)
);

AOI322xp5_ASAP7_75t_L g1027 ( 
.A1(n_1024),
.A2(n_907),
.A3(n_940),
.B1(n_970),
.B2(n_967),
.C1(n_973),
.C2(n_832),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1021),
.A2(n_941),
.B1(n_901),
.B2(n_970),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1020),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1022),
.B(n_975),
.Y(n_1030)
);

AOI322xp5_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_967),
.A3(n_873),
.B1(n_881),
.B2(n_844),
.C1(n_943),
.C2(n_937),
.Y(n_1031)
);

AOI21xp33_ASAP7_75t_SL g1032 ( 
.A1(n_1025),
.A2(n_816),
.B(n_910),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_1019),
.A2(n_826),
.B1(n_910),
.B2(n_856),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1030),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_1029),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1028),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1032),
.B(n_976),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1033),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1027),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

BUFx8_ASAP7_75t_SL g1041 ( 
.A(n_1029),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1029),
.Y(n_1042)
);

BUFx4_ASAP7_75t_SL g1043 ( 
.A(n_1029),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1030),
.Y(n_1044)
);

NAND4xp25_ASAP7_75t_L g1045 ( 
.A(n_1035),
.B(n_1026),
.C(n_810),
.D(n_976),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1035),
.B(n_947),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1041),
.B(n_828),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_1042),
.B(n_817),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_810),
.C(n_839),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_1034),
.B(n_811),
.C(n_865),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_1044),
.B(n_845),
.C(n_850),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1038),
.B(n_839),
.C(n_861),
.Y(n_1052)
);

AOI211x1_ASAP7_75t_L g1053 ( 
.A1(n_1037),
.A2(n_1043),
.B(n_1040),
.C(n_1036),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1043),
.B(n_882),
.C(n_889),
.Y(n_1054)
);

NOR4xp25_ASAP7_75t_L g1055 ( 
.A(n_1035),
.B(n_946),
.C(n_945),
.D(n_954),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1047),
.A2(n_1048),
.B(n_1046),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_L g1057 ( 
.A(n_1045),
.B(n_882),
.C(n_894),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_1052),
.B(n_882),
.C(n_883),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_1050),
.B(n_945),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1049),
.B(n_882),
.C(n_815),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1053),
.A2(n_923),
.B1(n_954),
.B2(n_884),
.C(n_947),
.Y(n_1061)
);

AND2x2_ASAP7_75t_SL g1062 ( 
.A(n_1054),
.B(n_824),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_1051),
.A2(n_923),
.B(n_912),
.Y(n_1063)
);

NOR2x1p5_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_1055),
.Y(n_1064)
);

NOR5xp2_ASAP7_75t_L g1065 ( 
.A(n_1063),
.B(n_946),
.C(n_909),
.D(n_916),
.E(n_915),
.Y(n_1065)
);

NAND5xp2_ASAP7_75t_L g1066 ( 
.A(n_1061),
.B(n_853),
.C(n_881),
.D(n_898),
.E(n_899),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_877),
.C(n_818),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_1058),
.A2(n_947),
.B(n_934),
.Y(n_1068)
);

NAND4xp75_ASAP7_75t_L g1069 ( 
.A(n_1062),
.B(n_897),
.C(n_898),
.D(n_899),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_SL g1070 ( 
.A1(n_1060),
.A2(n_908),
.B1(n_902),
.B2(n_931),
.C(n_955),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_L g1071 ( 
.A(n_1059),
.B(n_824),
.Y(n_1071)
);

AOI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1056),
.A2(n_932),
.B(n_824),
.C(n_884),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_1064),
.B(n_893),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1071),
.B(n_955),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1068),
.B(n_859),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1067),
.B(n_934),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1069),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_1072),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_939),
.B(n_896),
.Y(n_1079)
);

NOR2x1_ASAP7_75t_L g1080 ( 
.A(n_1066),
.B(n_931),
.Y(n_1080)
);

OAI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1065),
.A2(n_908),
.B1(n_819),
.B2(n_902),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1064),
.B(n_859),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_1073),
.Y(n_1083)
);

NAND4xp25_ASAP7_75t_SL g1084 ( 
.A(n_1082),
.B(n_939),
.C(n_903),
.D(n_904),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1075),
.A2(n_1074),
.B1(n_1079),
.B2(n_1081),
.C(n_1080),
.Y(n_1085)
);

AND3x4_ASAP7_75t_L g1086 ( 
.A(n_1076),
.B(n_934),
.C(n_892),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_SL g1087 ( 
.A(n_1073),
.B(n_956),
.C(n_951),
.Y(n_1087)
);

NOR2x1_ASAP7_75t_L g1088 ( 
.A(n_1082),
.B(n_893),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1078),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1082),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1082),
.Y(n_1091)
);

AO22x1_ASAP7_75t_SL g1092 ( 
.A1(n_1077),
.A2(n_884),
.B1(n_885),
.B2(n_880),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1089),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1083),
.A2(n_819),
.B1(n_902),
.B2(n_893),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1086),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1090),
.A2(n_902),
.B1(n_893),
.B2(n_951),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1091),
.Y(n_1097)
);

NAND4xp75_ASAP7_75t_L g1098 ( 
.A(n_1088),
.B(n_1085),
.C(n_1092),
.D(n_1084),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1095),
.A2(n_1087),
.B1(n_902),
.B2(n_956),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_1093),
.A2(n_885),
.B1(n_880),
.B2(n_886),
.Y(n_1100)
);

OA22x2_ASAP7_75t_L g1101 ( 
.A1(n_1097),
.A2(n_902),
.B1(n_880),
.B2(n_914),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1098),
.A2(n_896),
.B1(n_885),
.B2(n_897),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_1094),
.A2(n_886),
.B1(n_877),
.B2(n_897),
.Y(n_1103)
);

OA22x2_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1096),
.B1(n_877),
.B2(n_875),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1101),
.B(n_886),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1100),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_1105),
.A2(n_1099),
.B(n_1102),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1107),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1104),
.Y(n_1109)
);

AOI22x1_ASAP7_75t_L g1110 ( 
.A1(n_1109),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_1110)
);

OA22x2_ASAP7_75t_L g1111 ( 
.A1(n_1109),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1111),
.A2(n_878),
.B(n_897),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_161),
.B(n_164),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1113),
.B(n_886),
.Y(n_1114)
);

XOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_1112),
.B(n_165),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.C(n_175),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_1114),
.B(n_179),
.C(n_180),
.Y(n_1117)
);


endmodule