module fake_jpeg_6728_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_17),
.B1(n_22),
.B2(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_16),
.B1(n_22),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_16),
.B1(n_22),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_17),
.B1(n_25),
.B2(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_59),
.B1(n_39),
.B2(n_35),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_28),
.B1(n_15),
.B2(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_28),
.B1(n_15),
.B2(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_34),
.C(n_58),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_38),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_74),
.Y(n_100)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_78),
.B1(n_51),
.B2(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_33),
.B1(n_38),
.B2(n_15),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_19),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_97),
.B1(n_77),
.B2(n_74),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_51),
.A3(n_45),
.B1(n_60),
.B2(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_19),
.B(n_49),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_103),
.C(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_19),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_19),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_72),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_43),
.B1(n_28),
.B2(n_37),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_68),
.B1(n_67),
.B2(n_24),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_24),
.B(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_61),
.B1(n_75),
.B2(n_69),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_124),
.C(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_122),
.B1(n_123),
.B2(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_119),
.B(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_47),
.B1(n_37),
.B2(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_130),
.Y(n_149)
);

NAND2x1_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_138),
.Y(n_154)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_85),
.B1(n_99),
.B2(n_103),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_90),
.B1(n_83),
.B2(n_86),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_124),
.B1(n_122),
.B2(n_120),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_83),
.C(n_13),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_101),
.B(n_98),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_106),
.C(n_117),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_156),
.B1(n_101),
.B2(n_21),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.C(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_118),
.C(n_109),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_117),
.B1(n_105),
.B2(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_37),
.C(n_32),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_32),
.C(n_30),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_142),
.C(n_132),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_140),
.B(n_138),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_158),
.B(n_3),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_169),
.C(n_157),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_130),
.B1(n_126),
.B2(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_167),
.B1(n_165),
.B2(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_141),
.C(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_127),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_128),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_127),
.B(n_128),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_156),
.B(n_148),
.C(n_155),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_30),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_30),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_162),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_13),
.C(n_3),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_152),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_191),
.B(n_168),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_147),
.C(n_155),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_174),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.C(n_199),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_187),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_198),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_158),
.B(n_47),
.C(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_2),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.C(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_208),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_179),
.C(n_6),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_198),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_6),
.C(n_7),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_193),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_214),
.B(n_216),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_221),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_8),
.B(n_10),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_7),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_8),
.B(n_12),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_212),
.B(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_223),
.B(n_12),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_228),
.Y(n_230)
);


endmodule