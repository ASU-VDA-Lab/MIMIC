module fake_jpeg_9553_n_296 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_65)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_22),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_26),
.B1(n_22),
.B2(n_32),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_27),
.B1(n_34),
.B2(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_33),
.B1(n_23),
.B2(n_19),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_28),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_42),
.C(n_36),
.Y(n_101)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_70),
.Y(n_106)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_74),
.Y(n_115)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_41),
.B1(n_56),
.B2(n_21),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_40),
.B1(n_41),
.B2(n_23),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_19),
.B1(n_40),
.B2(n_27),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NOR4xp25_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_103),
.Y(n_116)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_42),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_28),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_60),
.B1(n_56),
.B2(n_44),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_56),
.B1(n_42),
.B2(n_41),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_78),
.B1(n_88),
.B2(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_28),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_123),
.B1(n_116),
.B2(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_145),
.B1(n_153),
.B2(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_137),
.B(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_89),
.B1(n_93),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_154),
.B1(n_133),
.B2(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_78),
.B1(n_102),
.B2(n_83),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_87),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_3),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_96),
.B1(n_103),
.B2(n_104),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_104),
.B1(n_70),
.B2(n_72),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_73),
.B1(n_36),
.B2(n_95),
.Y(n_154)
);

OR2x4_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_81),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_114),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_24),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_36),
.B1(n_24),
.B2(n_18),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_31),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_122),
.B(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_114),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_36),
.B(n_18),
.C(n_31),
.D(n_5),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_1),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_121),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_31),
.B(n_128),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_185),
.B1(n_158),
.B2(n_157),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_118),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_182),
.C(n_3),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_155),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_171),
.B(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_106),
.B1(n_129),
.B2(n_128),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_134),
.B1(n_162),
.B2(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_106),
.C(n_109),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_126),
.B1(n_112),
.B2(n_18),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_31),
.B(n_126),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_112),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_31),
.B(n_3),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_7),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_7),
.B(n_8),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_4),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_216),
.B1(n_169),
.B2(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_205),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_137),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_173),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_134),
.B1(n_4),
.B2(n_5),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_166),
.C(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_189),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_217),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_187),
.C(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_165),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_171),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_213),
.CI(n_185),
.CON(n_253),
.SN(n_253)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_179),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_209),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_180),
.B(n_174),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_193),
.B1(n_164),
.B2(n_172),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_207),
.B1(n_195),
.B2(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_205),
.B(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_245),
.B1(n_167),
.B2(n_172),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_244),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_232),
.Y(n_244)
);

OAI321xp33_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_216),
.A3(n_210),
.B1(n_208),
.B2(n_204),
.C(n_207),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_222),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_201),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_251),
.B(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_230),
.C(n_228),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.C(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_258),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_236),
.C(n_223),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_233),
.C(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_221),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_181),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_183),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_266),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_249),
.B(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

OAI221xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_262),
.B1(n_260),
.B2(n_263),
.C(n_15),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_249),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_275),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_196),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_240),
.C(n_10),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_8),
.Y(n_279)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_240),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_283),
.B1(n_10),
.B2(n_11),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_263),
.B1(n_11),
.B2(n_14),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_267),
.B(n_272),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_288),
.C(n_11),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_273),
.C(n_280),
.Y(n_288)
);

AOI211xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_290),
.B(n_286),
.C(n_288),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_15),
.B(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.Y(n_296)
);


endmodule