module fake_jpeg_1857_n_560 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_560);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_560;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_17),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_100),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_76),
.Y(n_124)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_30),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_98),
.Y(n_164)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_50),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_104),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_22),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_43),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_1),
.Y(n_148)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_52),
.B1(n_51),
.B2(n_22),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_106),
.A2(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_40),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_85),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_21),
.B1(n_36),
.B2(n_42),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_116),
.A2(n_140),
.B1(n_146),
.B2(n_78),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_52),
.B1(n_49),
.B2(n_38),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_131),
.B1(n_133),
.B2(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_54),
.A2(n_49),
.B1(n_28),
.B2(n_34),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_58),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_21),
.B1(n_36),
.B2(n_42),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_21),
.B(n_36),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_79),
.B(n_104),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_68),
.A2(n_41),
.B1(n_34),
.B2(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_141),
.B1(n_143),
.B2(n_165),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_53),
.A2(n_45),
.B1(n_44),
.B2(n_38),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_101),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_81),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_156),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_64),
.B(n_39),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_90),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_56),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_177),
.Y(n_234)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_170),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_181),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_94),
.B1(n_71),
.B2(n_72),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_119),
.B(n_107),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_183),
.B(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_152),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_189),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_135),
.B1(n_146),
.B2(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_196),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_105),
.B1(n_57),
.B2(n_95),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_152),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_116),
.A2(n_98),
.B1(n_114),
.B2(n_115),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_199),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_192),
.B(n_216),
.Y(n_277)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_83),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_194),
.B(n_214),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_125),
.A2(n_76),
.B1(n_73),
.B2(n_61),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_2),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_3),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_3),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_112),
.A2(n_142),
.B1(n_155),
.B2(n_108),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_222),
.B1(n_229),
.B2(n_166),
.Y(n_275)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_3),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_215),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_124),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_123),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_226),
.Y(n_262)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_160),
.A2(n_24),
.B1(n_5),
.B2(n_7),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_161),
.B1(n_129),
.B2(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_230),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_145),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_154),
.A2(n_24),
.B1(n_5),
.B2(n_8),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_154),
.B(n_4),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_174),
.B1(n_178),
.B2(n_194),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_168),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g318 ( 
.A1(n_239),
.A2(n_201),
.B(n_172),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_192),
.A2(n_126),
.B1(n_168),
.B2(n_129),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_181),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_173),
.A2(n_166),
.B1(n_123),
.B2(n_145),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_194),
.B1(n_224),
.B2(n_171),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_123),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_280),
.C(n_201),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_175),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_214),
.B1(n_184),
.B2(n_189),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_180),
.B(n_191),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_200),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_282),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_219),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_291),
.Y(n_356)
);

AO21x2_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_238),
.B(n_241),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_180),
.B1(n_173),
.B2(n_214),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_297),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_298),
.A2(n_311),
.B1(n_313),
.B2(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_173),
.B(n_223),
.C(n_193),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_300),
.A2(n_272),
.B(n_278),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_227),
.B1(n_217),
.B2(n_207),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_236),
.Y(n_343)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_222),
.B1(n_179),
.B2(n_188),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_303),
.A2(n_308),
.B1(n_326),
.B2(n_237),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_255),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_304),
.B(n_307),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_245),
.B1(n_258),
.B2(n_274),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_239),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_309),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_262),
.A2(n_197),
.B1(n_220),
.B2(n_226),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_218),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_243),
.A2(n_198),
.B1(n_213),
.B2(n_24),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_312),
.B(n_314),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_255),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_267),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_319),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_263),
.B(n_233),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_320),
.B(n_321),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_232),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_323),
.Y(n_339)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_172),
.C(n_10),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_331),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_234),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_327),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_232),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_328),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_12),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_330),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_13),
.C(n_14),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_333),
.Y(n_350)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_258),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_263),
.C(n_251),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_335),
.B(n_332),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_336),
.A2(n_334),
.B1(n_240),
.B2(n_273),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_340),
.A2(n_345),
.B(n_355),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_247),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_372),
.C(n_288),
.Y(n_379)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_360),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_293),
.A2(n_245),
.B(n_284),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_289),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_366),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_246),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_363),
.A2(n_374),
.B(n_305),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_368),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_290),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_292),
.A2(n_273),
.B1(n_240),
.B2(n_268),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_259),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_300),
.A2(n_272),
.B(n_237),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_306),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_373),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_403),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_311),
.B1(n_306),
.B2(n_305),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_387),
.B1(n_401),
.B2(n_409),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_391),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_372),
.C(n_342),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_386),
.C(n_397),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_355),
.B(n_340),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_385),
.A2(n_395),
.B(n_412),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_288),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_327),
.B1(n_325),
.B2(n_313),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_331),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_399),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_390),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_346),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_364),
.A2(n_308),
.B1(n_330),
.B2(n_291),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_350),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_394),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_350),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_302),
.B(n_285),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_361),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_396),
.B(n_400),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_333),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_335),
.B(n_323),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_360),
.B(n_326),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_336),
.A2(n_316),
.B1(n_286),
.B2(n_310),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_406),
.B1(n_410),
.B2(n_414),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_337),
.B(n_321),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_404),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_320),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_411),
.C(n_338),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_351),
.A2(n_294),
.B1(n_315),
.B2(n_236),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_249),
.Y(n_407)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_352),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_336),
.A2(n_249),
.B1(n_231),
.B2(n_297),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_13),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_371),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_15),
.Y(n_413)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_365),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g418 ( 
.A(n_403),
.B(n_347),
.CI(n_351),
.CON(n_418),
.SN(n_418)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_418),
.B(n_408),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_423),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_441),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_367),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_368),
.B1(n_359),
.B2(n_363),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_427),
.A2(n_428),
.B1(n_433),
.B2(n_443),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_393),
.A2(n_394),
.B1(n_392),
.B2(n_409),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_398),
.A2(n_374),
.B(n_345),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_431),
.B(n_391),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_398),
.A2(n_359),
.B(n_357),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_357),
.C(n_344),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_446),
.C(n_395),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_387),
.A2(n_339),
.B1(n_343),
.B2(n_356),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_386),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_439),
.Y(n_454)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_438),
.Y(n_450)
);

XNOR2x1_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_338),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_344),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_381),
.A2(n_356),
.B1(n_369),
.B2(n_362),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_392),
.A2(n_369),
.B1(n_362),
.B2(n_377),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_445),
.A2(n_402),
.B1(n_410),
.B2(n_412),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_371),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_452),
.A2(n_465),
.B1(n_466),
.B2(n_469),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_444),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_453),
.B(n_468),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_464),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_417),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_457),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_411),
.C(n_396),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_471),
.C(n_451),
.Y(n_482)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_390),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_463),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_441),
.B(n_389),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_428),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_425),
.A2(n_408),
.B1(n_406),
.B2(n_404),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_467),
.B(n_418),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_442),
.B(n_400),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_429),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_470),
.A2(n_430),
.B(n_434),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_432),
.C(n_435),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_472),
.A2(n_473),
.B1(n_427),
.B2(n_431),
.Y(n_480)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_437),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_474),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_479),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_420),
.Y(n_479)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_485),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_484),
.A2(n_495),
.B(n_497),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_421),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_416),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_458),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_416),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_475),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_448),
.A2(n_434),
.B1(n_419),
.B2(n_418),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_488),
.A2(n_484),
.B1(n_490),
.B2(n_495),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_SL g489 ( 
.A(n_457),
.B(n_467),
.C(n_456),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_491),
.C(n_454),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_446),
.C(n_439),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_448),
.A2(n_419),
.B1(n_407),
.B2(n_413),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_492),
.A2(n_465),
.B1(n_452),
.B2(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_493),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_414),
.B(n_377),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_457),
.A2(n_370),
.B(n_17),
.Y(n_497)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_496),
.Y(n_503)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_503),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_509),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_481),
.A2(n_464),
.B1(n_455),
.B2(n_473),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_505),
.A2(n_510),
.B1(n_513),
.B2(n_491),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_454),
.C(n_466),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_482),
.C(n_489),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_449),
.B1(n_450),
.B2(n_474),
.Y(n_508)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_508),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_481),
.A2(n_370),
.B(n_17),
.C(n_18),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_494),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_16),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_511),
.Y(n_520)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_487),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_515),
.A2(n_476),
.B1(n_485),
.B2(n_513),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_515),
.B(n_493),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_525),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_517),
.B(n_500),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_498),
.A2(n_490),
.B(n_483),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_522),
.A2(n_523),
.B(n_512),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_498),
.A2(n_488),
.B(n_497),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_516),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_501),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_511),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_529),
.B(n_530),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_499),
.C(n_514),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_531),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_502),
.C(n_499),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_533),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_504),
.C(n_506),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_534),
.A2(n_538),
.B(n_541),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_528),
.B(n_505),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_522),
.C(n_518),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_519),
.B(n_503),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_537),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_500),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_547),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_530),
.C(n_526),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_532),
.B(n_524),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_540),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_544),
.B(n_531),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_551),
.Y(n_553)
);

AOI21xp33_ASAP7_75t_L g551 ( 
.A1(n_543),
.A2(n_518),
.B(n_523),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_552),
.B(n_542),
.C(n_546),
.Y(n_554)
);

AOI31xp67_ASAP7_75t_L g556 ( 
.A1(n_554),
.A2(n_535),
.A3(n_534),
.B(n_525),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_553),
.A2(n_550),
.B(n_546),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_555),
.B(n_556),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_520),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_558),
.B(n_520),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_512),
.B(n_509),
.Y(n_560)
);


endmodule