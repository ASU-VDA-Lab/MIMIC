module fake_jpeg_13214_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g160 ( 
.A(n_54),
.Y(n_160)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_20),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_105),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_29),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_111),
.Y(n_158)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_113),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_20),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_23),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_155),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_105),
.A2(n_38),
.B(n_50),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_150),
.B(n_16),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_59),
.A2(n_43),
.B1(n_38),
.B2(n_50),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_173),
.B1(n_175),
.B2(n_179),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_108),
.A2(n_52),
.B1(n_50),
.B2(n_38),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_24),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_178),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_79),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_56),
.A2(n_51),
.B1(n_26),
.B2(n_31),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_42),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_95),
.A2(n_35),
.B1(n_31),
.B2(n_51),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_47),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_183),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_60),
.A2(n_35),
.B1(n_45),
.B2(n_25),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_81),
.B1(n_103),
.B2(n_106),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_98),
.B(n_25),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_184),
.Y(n_281)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_122),
.A2(n_24),
.B1(n_45),
.B2(n_74),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_122),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_193),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_119),
.B(n_0),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_202),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_218),
.Y(n_265)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_198),
.Y(n_299)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_200),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_0),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_203),
.B(n_211),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_206),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_136),
.Y(n_207)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_213),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_132),
.B(n_178),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_113),
.B1(n_104),
.B2(n_102),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_212),
.A2(n_214),
.B1(n_236),
.B2(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_110),
.B1(n_39),
.B2(n_84),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_221),
.A2(n_124),
.B1(n_170),
.B2(n_156),
.Y(n_270)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_226),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_1),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_128),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_227),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_140),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_163),
.B(n_2),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_159),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_151),
.B1(n_131),
.B2(n_115),
.Y(n_278)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_232),
.Y(n_286)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_234),
.Y(n_291)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_172),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_175),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_114),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_160),
.B(n_2),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_152),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_130),
.C(n_8),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_6),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_6),
.Y(n_274)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_129),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_245),
.Y(n_284)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_149),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_246),
.Y(n_295)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_6),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_172),
.B(n_160),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_274),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_191),
.A2(n_145),
.B1(n_118),
.B2(n_117),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_261),
.A2(n_209),
.B(n_246),
.C(n_244),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_272),
.B1(n_277),
.B2(n_280),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_177),
.B1(n_166),
.B2(n_157),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_201),
.A2(n_177),
.B1(n_166),
.B2(n_157),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_189),
.B1(n_200),
.B2(n_232),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_227),
.B(n_7),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_297),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_186),
.A2(n_151),
.B1(n_167),
.B2(n_130),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_198),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_225),
.B(n_7),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_247),
.C(n_245),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_7),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_271),
.A2(n_243),
.B1(n_230),
.B2(n_195),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_221),
.B1(n_242),
.B2(n_202),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_340),
.B1(n_283),
.B2(n_295),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_305),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_196),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_194),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_226),
.B(n_215),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_308),
.A2(n_332),
.B(n_252),
.Y(n_364)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_298),
.B(n_274),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_311),
.A2(n_313),
.B(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_314),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_205),
.B(n_222),
.C(n_188),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_234),
.Y(n_314)
);

XOR2x2_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_207),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_339),
.C(n_316),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_333),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_318),
.B(n_326),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_322),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_273),
.B(n_218),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_193),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_192),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_324),
.Y(n_349)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_253),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_325),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_297),
.B(n_185),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_328),
.Y(n_354)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_254),
.B(n_199),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_329),
.B(n_331),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_251),
.B(n_217),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_270),
.A2(n_208),
.B(n_235),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_250),
.B1(n_264),
.B2(n_284),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_335),
.B(n_337),
.Y(n_345)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_338),
.B(n_341),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_223),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_265),
.A2(n_204),
.B1(n_8),
.B2(n_9),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_353),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_302),
.A2(n_300),
.B1(n_320),
.B2(n_315),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_300),
.A2(n_261),
.B1(n_267),
.B2(n_265),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_259),
.C(n_261),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_367),
.C(n_372),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_261),
.B1(n_259),
.B2(n_281),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_268),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_359),
.A2(n_364),
.B(n_366),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_286),
.B1(n_281),
.B2(n_269),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_360),
.A2(n_365),
.B1(n_330),
.B2(n_262),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_323),
.A2(n_250),
.B1(n_288),
.B2(n_284),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_306),
.A2(n_319),
.B1(n_322),
.B2(n_327),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_257),
.C(n_275),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_317),
.B1(n_313),
.B2(n_337),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_306),
.A2(n_291),
.B(n_299),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g398 ( 
.A1(n_370),
.A2(n_371),
.B(n_290),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_306),
.A2(n_288),
.B(n_266),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_266),
.C(n_276),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_341),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_264),
.B1(n_252),
.B2(n_268),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_374),
.A2(n_328),
.B1(n_336),
.B2(n_317),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_294),
.C(n_262),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_9),
.C(n_11),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_381),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_355),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_360),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_384),
.A2(n_386),
.B(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_303),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_392),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_357),
.A2(n_308),
.B(n_317),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_317),
.B1(n_324),
.B2(n_309),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_387),
.A2(n_388),
.B1(n_405),
.B2(n_411),
.Y(n_429)
);

OA22x2_ASAP7_75t_L g444 ( 
.A1(n_389),
.A2(n_374),
.B1(n_368),
.B2(n_365),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_354),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_390),
.B(n_396),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_413),
.C(n_372),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_338),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_333),
.B(n_307),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_366),
.A2(n_312),
.B(n_310),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_395),
.A2(n_398),
.B(n_349),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_276),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_362),
.B(n_287),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_397),
.B(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_401),
.Y(n_417)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_287),
.Y(n_403)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_404),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_350),
.A2(n_290),
.B1(n_294),
.B2(n_287),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_407),
.Y(n_432)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_7),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_410),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_8),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_359),
.A2(n_294),
.B1(n_11),
.B2(n_12),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_349),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_379),
.A2(n_344),
.B1(n_373),
.B2(n_356),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_426),
.B1(n_437),
.B2(n_446),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_397),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_424),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_405),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_385),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_379),
.A2(n_346),
.B1(n_359),
.B2(n_371),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_400),
.A2(n_347),
.B1(n_353),
.B2(n_368),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_398),
.B1(n_401),
.B2(n_394),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_383),
.A2(n_376),
.B(n_368),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_396),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_438),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_345),
.C(n_372),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_443),
.C(n_367),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_369),
.B1(n_346),
.B2(n_368),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_403),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_393),
.B(n_378),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_343),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_392),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_442),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_384),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_345),
.C(n_378),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_387),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_383),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_412),
.A2(n_370),
.B1(n_377),
.B2(n_367),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_449),
.A2(n_450),
.B1(n_388),
.B2(n_444),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_475),
.Y(n_484)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_454),
.A2(n_459),
.B1(n_468),
.B2(n_422),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_466),
.C(n_471),
.Y(n_478)
);

OAI322xp33_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_409),
.A3(n_408),
.B1(n_407),
.B2(n_406),
.C1(n_399),
.C2(n_402),
.Y(n_458)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_458),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_414),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_439),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_464),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_384),
.C(n_395),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_348),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_467),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_398),
.B1(n_381),
.B2(n_380),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_417),
.A2(n_421),
.B1(n_437),
.B2(n_426),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_469),
.A2(n_428),
.B1(n_442),
.B2(n_430),
.Y(n_481)
);

BUFx12_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_470),
.Y(n_497)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_472),
.A2(n_473),
.B1(n_436),
.B2(n_410),
.Y(n_499)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_425),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_474),
.Y(n_498)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_451),
.A2(n_429),
.B1(n_417),
.B2(n_441),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_477),
.A2(n_481),
.B1(n_495),
.B2(n_473),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_440),
.C(n_423),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_483),
.C(n_488),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_420),
.C(n_438),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_450),
.A2(n_420),
.B1(n_415),
.B2(n_418),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_487),
.A2(n_489),
.B1(n_493),
.B2(n_464),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_419),
.C(n_415),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_466),
.B(n_445),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_490),
.B(n_494),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_450),
.A2(n_418),
.B1(n_434),
.B2(n_444),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_436),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_386),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_469),
.A2(n_447),
.B1(n_472),
.B2(n_453),
.Y(n_495)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_447),
.C(n_455),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_501),
.B(n_503),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_455),
.C(n_461),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_462),
.C(n_460),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_508),
.C(n_511),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_492),
.Y(n_505)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_460),
.Y(n_506)
);

XNOR2x1_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_509),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_484),
.C(n_490),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_487),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_510),
.B(n_517),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_465),
.C(n_456),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_482),
.A2(n_448),
.B(n_451),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_512),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_444),
.Y(n_513)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_515),
.B(n_496),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_493),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_495),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_482),
.B1(n_500),
.B2(n_486),
.Y(n_522)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_519),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_531),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_532),
.Y(n_540)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_514),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_529),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_497),
.C(n_479),
.Y(n_529)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_534),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_507),
.A2(n_479),
.B1(n_489),
.B2(n_416),
.Y(n_531)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_504),
.Y(n_534)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_503),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_521),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_527),
.A2(n_498),
.B1(n_513),
.B2(n_508),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_545),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_525),
.A2(n_502),
.B(n_515),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_542),
.A2(n_550),
.B(n_363),
.Y(n_558)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_502),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_546),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_513),
.C(n_439),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_535),
.B(n_470),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_470),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_547),
.B(n_548),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_529),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_533),
.Y(n_549)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_549),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_382),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_531),
.C(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_556),
.Y(n_564)
);

AO22x1_ASAP7_75t_L g554 ( 
.A1(n_539),
.A2(n_520),
.B1(n_524),
.B2(n_411),
.Y(n_554)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_554),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_363),
.C(n_348),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_558),
.B(n_546),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_537),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_560),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_16),
.C(n_12),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_552),
.B(n_549),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_552),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_563),
.B(n_566),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_538),
.C(n_540),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_568),
.B(n_551),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_570),
.B(n_571),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_564),
.A2(n_561),
.B(n_557),
.Y(n_572)
);

NAND4xp25_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_567),
.C(n_565),
.D(n_551),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_574),
.A2(n_569),
.B(n_553),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_573),
.B(n_547),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_560),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_577),
.A2(n_554),
.B(n_559),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_12),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_14),
.C(n_573),
.Y(n_580)
);


endmodule