module fake_jpeg_1095_n_676 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_676);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_676;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_57),
.C(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_59),
.B(n_63),
.Y(n_155)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g179 ( 
.A(n_65),
.Y(n_179)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_70),
.Y(n_200)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_72),
.Y(n_206)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g162 ( 
.A(n_80),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_81),
.B(n_87),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_10),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_90),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_91),
.B(n_117),
.Y(n_158)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_94),
.Y(n_137)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_98),
.Y(n_227)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_33),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_104),
.Y(n_226)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_107),
.Y(n_230)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_123),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_113),
.B(n_0),
.Y(n_229)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_21),
.B(n_10),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx5_ASAP7_75t_SL g193 ( 
.A(n_119),
.Y(n_193)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_48),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_25),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_130),
.B(n_131),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g131 ( 
.A(n_37),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_57),
.B1(n_24),
.B2(n_25),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_132),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_134),
.B(n_154),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_37),
.B1(n_53),
.B2(n_56),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_135),
.B(n_111),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_37),
.B1(n_31),
.B2(n_22),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_22),
.B1(n_55),
.B2(n_56),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_68),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_50),
.B1(n_40),
.B2(n_36),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_145),
.A2(n_149),
.B1(n_183),
.B2(n_196),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_40),
.B1(n_36),
.B2(n_27),
.Y(n_149)
);

AND2x4_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_0),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_152),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_27),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_81),
.B(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_161),
.B(n_169),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_172),
.A2(n_4),
.B1(n_141),
.B2(n_143),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_10),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_178),
.B(n_180),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_11),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_62),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_72),
.B(n_19),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_60),
.A2(n_8),
.B1(n_18),
.B2(n_16),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_189),
.A2(n_207),
.B1(n_216),
.B2(n_166),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_58),
.B(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_192),
.B(n_222),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_62),
.A2(n_125),
.B1(n_77),
.B2(n_131),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_8),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_93),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_199),
.B(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_79),
.B(n_19),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_61),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_82),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_215),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_125),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_209),
.A2(n_214),
.B1(n_1),
.B2(n_3),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_83),
.A2(n_5),
.B1(n_13),
.B2(n_12),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_84),
.B(n_15),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_64),
.A2(n_5),
.B1(n_12),
.B2(n_15),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_88),
.B(n_5),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_98),
.B(n_0),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_228),
.B(n_4),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_137),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_268),
.Y(n_322)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_234),
.Y(n_351)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g325 ( 
.A(n_236),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_238),
.Y(n_339)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_241),
.Y(n_348)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_179),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_244),
.B(n_251),
.C(n_275),
.Y(n_371)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_245),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_246),
.Y(n_361)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_247),
.Y(n_356)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_152),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_250),
.B(n_259),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_155),
.B(n_1),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_252),
.B(n_272),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_254),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_255),
.Y(n_362)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_138),
.Y(n_256)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_152),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_139),
.Y(n_260)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_260),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_207),
.A2(n_109),
.B1(n_107),
.B2(n_104),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_261),
.Y(n_363)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_262),
.Y(n_358)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_264),
.Y(n_360)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_156),
.Y(n_265)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_265),
.Y(n_364)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_266),
.Y(n_377)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_267),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_158),
.A2(n_80),
.B(n_65),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_271),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_144),
.B(n_1),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_162),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_273),
.B(n_291),
.Y(n_359)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_274),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_179),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_186),
.A2(n_3),
.B(n_4),
.C(n_151),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_298),
.B(n_300),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_185),
.B(n_3),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_279),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_150),
.B(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_294),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_284),
.B(n_290),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_189),
.A2(n_4),
.B1(n_204),
.B2(n_160),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_285),
.A2(n_295),
.B1(n_297),
.B2(n_299),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_289),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_288),
.Y(n_326)
);

BUFx4f_ASAP7_75t_SL g289 ( 
.A(n_160),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_133),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_175),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_292),
.A2(n_309),
.B1(n_310),
.B2(n_313),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_185),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_293),
.B(n_296),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_135),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_200),
.A2(n_225),
.B1(n_153),
.B2(n_147),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_176),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_168),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_170),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_171),
.B(n_177),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_172),
.B(n_149),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_302),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_137),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_165),
.A2(n_166),
.B1(n_174),
.B2(n_173),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_303),
.A2(n_307),
.B1(n_311),
.B2(n_314),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_195),
.B(n_221),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_305),
.Y(n_338)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_217),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_308),
.Y(n_378)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_148),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_168),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_157),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_147),
.B(n_153),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_317),
.Y(n_329)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_148),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_200),
.A2(n_206),
.B1(n_217),
.B2(n_221),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_140),
.A2(n_145),
.B(n_209),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_187),
.C(n_193),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_165),
.B(n_174),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_284),
.A2(n_214),
.B1(n_173),
.B2(n_157),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_319),
.A2(n_323),
.B1(n_374),
.B2(n_289),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_163),
.B1(n_187),
.B2(n_183),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_279),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_164),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_354),
.C(n_370),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_163),
.B1(n_227),
.B2(n_142),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_352),
.B1(n_357),
.B2(n_367),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_231),
.A2(n_142),
.B1(n_194),
.B2(n_227),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_SL g354 ( 
.A(n_252),
.B(n_193),
.C(n_146),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_292),
.A2(n_224),
.B1(n_202),
.B2(n_226),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_233),
.A2(n_194),
.B1(n_181),
.B2(n_190),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_233),
.A2(n_181),
.B1(n_190),
.B2(n_202),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_376),
.B1(n_306),
.B2(n_311),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_253),
.B(n_224),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_232),
.A2(n_315),
.B1(n_239),
.B2(n_309),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_272),
.A2(n_226),
.B1(n_164),
.B2(n_146),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_341),
.B(n_280),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_380),
.B(n_386),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_263),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_399),
.C(n_418),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_331),
.A2(n_276),
.B(n_237),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_385),
.A2(n_391),
.B(n_428),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_359),
.B(n_283),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_322),
.B(n_374),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_387),
.A2(n_402),
.B(n_426),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_327),
.A2(n_281),
.B1(n_269),
.B2(n_317),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_389),
.A2(n_395),
.B1(n_363),
.B2(n_319),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_304),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_398),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_324),
.B(n_366),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_393),
.B(n_403),
.Y(n_445)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_330),
.B(n_241),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_396),
.B(n_243),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_323),
.A2(n_289),
.B1(n_246),
.B2(n_279),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_397),
.A2(n_405),
.B1(n_408),
.B2(n_415),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_329),
.B(n_248),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_329),
.B(n_258),
.C(n_262),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_268),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_400),
.Y(n_441)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_334),
.A2(n_312),
.B(n_249),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_278),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_337),
.A2(n_313),
.B1(n_308),
.B2(n_256),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_407),
.B(n_412),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_327),
.A2(n_299),
.B1(n_290),
.B2(n_265),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_360),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_410),
.Y(n_436)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_267),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_236),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_416),
.Y(n_448)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_324),
.B(n_312),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_371),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_420),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_235),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_236),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_419),
.Y(n_443)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_266),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_423),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_322),
.B(n_343),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_372),
.C(n_361),
.Y(n_434)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_270),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_428),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_238),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_425),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_322),
.A2(n_240),
.B(n_297),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_427),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_372),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_354),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_430),
.B(n_451),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_395),
.A2(n_337),
.B1(n_357),
.B2(n_363),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_431),
.A2(n_464),
.B1(n_405),
.B2(n_408),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_469),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_439),
.B1(n_452),
.B2(n_468),
.Y(n_473)
);

AOI32xp33_ASAP7_75t_L g438 ( 
.A1(n_400),
.A2(n_349),
.A3(n_361),
.B1(n_320),
.B2(n_326),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_438),
.B(n_459),
.C(n_385),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_394),
.B1(n_401),
.B2(n_387),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_318),
.C(n_349),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_442),
.B(n_450),
.C(n_457),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_373),
.C(n_368),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_382),
.B(n_376),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_392),
.A2(n_340),
.B1(n_345),
.B2(n_342),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_398),
.B(n_325),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_SL g459 ( 
.A(n_417),
.B(n_325),
.C(n_302),
.Y(n_459)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_245),
.C(n_365),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_365),
.C(n_350),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_391),
.A2(n_288),
.B1(n_247),
.B2(n_345),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_383),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_400),
.A2(n_274),
.B1(n_264),
.B2(n_242),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_350),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_471),
.A2(n_480),
.B1(n_485),
.B2(n_486),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_399),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_499),
.C(n_507),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_455),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_474),
.B(n_484),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_509),
.Y(n_512)
);

OAI32xp33_ASAP7_75t_L g477 ( 
.A1(n_433),
.A2(n_393),
.A3(n_391),
.B1(n_421),
.B2(n_411),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_479),
.Y(n_518)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_441),
.A2(n_400),
.B1(n_389),
.B2(n_402),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_483),
.A2(n_497),
.B(n_510),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_460),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_397),
.B1(n_400),
.B2(n_416),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_452),
.A2(n_426),
.B1(n_407),
.B2(n_412),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_444),
.B(n_420),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_487),
.B(n_445),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_437),
.A2(n_424),
.B1(n_409),
.B2(n_418),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_488),
.A2(n_492),
.B1(n_494),
.B2(n_504),
.Y(n_525)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_490),
.Y(n_526)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_433),
.A2(n_414),
.B1(n_406),
.B2(n_427),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_460),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_493),
.B(n_509),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_449),
.A2(n_410),
.B1(n_404),
.B2(n_381),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_498),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_325),
.B(n_423),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_432),
.B(n_332),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_332),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_434),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_404),
.Y(n_502)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_431),
.A2(n_328),
.B1(n_344),
.B2(n_356),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_447),
.A2(n_328),
.B1(n_344),
.B2(n_356),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_505),
.A2(n_504),
.B1(n_492),
.B2(n_494),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_441),
.A2(n_379),
.B1(n_377),
.B2(n_286),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_506),
.A2(n_466),
.B1(n_468),
.B2(n_464),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_450),
.B(n_255),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_310),
.C(n_377),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_457),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_462),
.B(n_362),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_465),
.A2(n_362),
.B(n_257),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_511),
.A2(n_527),
.B1(n_529),
.B2(n_530),
.Y(n_561)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_513),
.B(n_523),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_483),
.A2(n_453),
.B1(n_448),
.B2(n_429),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_517),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_520),
.B(n_489),
.Y(n_552)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_481),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_503),
.A2(n_451),
.B1(n_447),
.B2(n_453),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_473),
.A2(n_443),
.B1(n_458),
.B2(n_429),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_488),
.A2(n_443),
.B1(n_458),
.B2(n_438),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_533),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_442),
.B1(n_454),
.B2(n_463),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_534),
.A2(n_543),
.B1(n_511),
.B2(n_521),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_478),
.A2(n_469),
.B1(n_461),
.B2(n_463),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_480),
.A2(n_459),
.B1(n_435),
.B2(n_440),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_482),
.A2(n_435),
.B1(n_440),
.B2(n_277),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_497),
.A2(n_510),
.B(n_506),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_475),
.B(n_496),
.Y(n_553)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_542),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_499),
.B(n_507),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_547),
.Y(n_571)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_472),
.Y(n_545)
);

BUFx24_ASAP7_75t_SL g564 ( 
.A(n_545),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_502),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_489),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_562),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_552),
.B(n_556),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_475),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_554),
.B(n_572),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_515),
.Y(n_556)
);

FAx1_ASAP7_75t_SL g557 ( 
.A(n_517),
.B(n_495),
.CI(n_477),
.CON(n_557),
.SN(n_557)
);

AOI21xp33_ASAP7_75t_L g589 ( 
.A1(n_557),
.A2(n_575),
.B(n_539),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_495),
.C(n_501),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_560),
.C(n_567),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_529),
.A2(n_491),
.B1(n_498),
.B2(n_508),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_559),
.A2(n_563),
.B1(n_576),
.B2(n_525),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_532),
.C(n_534),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_519),
.B(n_527),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_512),
.Y(n_565)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_565),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_536),
.B(n_521),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_566),
.B(n_568),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_546),
.C(n_518),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_541),
.Y(n_568)
);

NAND2x1_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_540),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_569),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_535),
.Y(n_570)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_570),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_516),
.B(n_541),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_522),
.B(n_546),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_573),
.B(n_531),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_522),
.B(n_514),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_574),
.B(n_562),
.Y(n_603)
);

FAx1_ASAP7_75t_SL g575 ( 
.A(n_539),
.B(n_514),
.CI(n_547),
.CON(n_575),
.SN(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_531),
.A2(n_518),
.B1(n_526),
.B2(n_513),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_535),
.Y(n_577)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_577),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_520),
.B(n_538),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g596 ( 
.A(n_578),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_571),
.Y(n_580)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_581),
.B(n_603),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_555),
.Y(n_583)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_583),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_587),
.B(n_574),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_561),
.Y(n_588)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_589),
.A2(n_569),
.B(n_558),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_554),
.B(n_537),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_598),
.Y(n_605)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_594),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_549),
.A2(n_528),
.B1(n_553),
.B2(n_575),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_600),
.B1(n_557),
.B2(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_597),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_551),
.B(n_528),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_576),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_599),
.B(n_566),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_572),
.A2(n_568),
.B1(n_549),
.B2(n_573),
.Y(n_600)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_604),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_579),
.Y(n_606)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_559),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_607),
.B(n_610),
.Y(n_635)
);

MAJx2_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_613),
.C(n_605),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_560),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_596),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_611),
.B(n_617),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_SL g629 ( 
.A1(n_614),
.A2(n_623),
.B(n_586),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_585),
.B(n_551),
.C(n_550),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_593),
.C(n_598),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_593),
.C(n_582),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_581),
.A2(n_557),
.B1(n_570),
.B2(n_577),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_620),
.A2(n_616),
.B1(n_613),
.B2(n_609),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_603),
.B(n_564),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_612),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_592),
.Y(n_623)
);

BUFx24_ASAP7_75t_SL g624 ( 
.A(n_587),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_624),
.B(n_621),
.Y(n_639)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_623),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_637),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_615),
.A2(n_600),
.B1(n_590),
.B2(n_602),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_627),
.A2(n_632),
.B1(n_633),
.B2(n_626),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_628),
.B(n_630),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_629),
.B(n_640),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_617),
.B(n_582),
.C(n_586),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_630),
.B(n_631),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_619),
.B(n_601),
.C(n_602),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_618),
.A2(n_601),
.B1(n_620),
.B2(n_614),
.Y(n_632)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_606),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_638),
.B(n_641),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_639),
.B(n_628),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_616),
.A2(n_622),
.B(n_608),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_644),
.B(n_645),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_635),
.B(n_605),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_634),
.Y(n_646)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_646),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_641),
.B(n_625),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_648),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_649),
.A2(n_651),
.B(n_652),
.Y(n_656)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_650),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_632),
.A2(n_627),
.B(n_633),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_638),
.C(n_640),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_637),
.B(n_634),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_653),
.B(n_652),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_647),
.A2(n_643),
.B(n_642),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_657),
.Y(n_663)
);

INVxp33_ASAP7_75t_SL g658 ( 
.A(n_654),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_658),
.B(n_660),
.Y(n_666)
);

FAx1_ASAP7_75t_SL g664 ( 
.A(n_659),
.B(n_661),
.CI(n_658),
.CON(n_664),
.SN(n_664)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_664),
.B(n_665),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_656),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_662),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_667),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_666),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_670),
.A2(n_655),
.B(n_654),
.Y(n_671)
);

BUFx24_ASAP7_75t_SL g673 ( 
.A(n_671),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_669),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_672),
.B(n_663),
.C(n_668),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_674),
.A2(n_651),
.B(n_643),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_675),
.Y(n_676)
);


endmodule