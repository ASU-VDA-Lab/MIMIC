module fake_jpeg_18693_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_34),
.B1(n_25),
.B2(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_22),
.B1(n_32),
.B2(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_58),
.B1(n_64),
.B2(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_20),
.B1(n_28),
.B2(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_24),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_26),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_37),
.C(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_21),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_76),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_41),
.B1(n_20),
.B2(n_23),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_91),
.B1(n_100),
.B2(n_27),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_88),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_41),
.B(n_24),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_81),
.B(n_97),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_22),
.B1(n_18),
.B2(n_32),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_41),
.B1(n_31),
.B2(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_21),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_40),
.B1(n_23),
.B2(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_26),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_43),
.B(n_31),
.C(n_16),
.D(n_30),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_26),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_28),
.B1(n_37),
.B2(n_29),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_106),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_54),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_31),
.Y(n_124)
);

NAND2x1_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_43),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_30),
.B(n_17),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_47),
.B(n_53),
.C(n_29),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_110),
.A2(n_71),
.B(n_104),
.C(n_74),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_37),
.B1(n_55),
.B2(n_27),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_116),
.B1(n_132),
.B2(n_133),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_1),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_106),
.B1(n_107),
.B2(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_105),
.B1(n_75),
.B2(n_81),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_30),
.B1(n_17),
.B2(n_16),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_91),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_162),
.B1(n_166),
.B2(n_121),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_108),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_145),
.B(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_112),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_100),
.B(n_68),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_84),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_151),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_112),
.B(n_115),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_156),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_12),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_159),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_68),
.B(n_2),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_17),
.B(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_114),
.B(n_120),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_94),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_1),
.B(n_69),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_70),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_126),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_136),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_90),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_129),
.B1(n_124),
.B2(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_4),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_124),
.B(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_163),
.B1(n_160),
.B2(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_127),
.Y(n_220)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_136),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_156),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_135),
.B1(n_121),
.B2(n_114),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_139),
.B1(n_169),
.B2(n_159),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_130),
.B(n_119),
.Y(n_193)
);

AOI22x1_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_127),
.B1(n_7),
.B2(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_119),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_146),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_11),
.B(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_90),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_209),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_210),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_191),
.A2(n_139),
.B1(n_140),
.B2(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_143),
.C(n_154),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_153),
.B1(n_158),
.B2(n_142),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_212),
.B1(n_193),
.B2(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_153),
.B1(n_167),
.B2(n_162),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_153),
.C(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_127),
.C(n_7),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_6),
.C(n_10),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_227),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_11),
.B(n_14),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_226),
.B(n_188),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_171),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_188),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_214),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_186),
.B(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_244),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_218),
.B1(n_193),
.B2(n_189),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_219),
.B1(n_216),
.B2(n_175),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_246),
.A2(n_181),
.B1(n_183),
.B2(n_206),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_175),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_181),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_250),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_209),
.C(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_252),
.C(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_208),
.C(n_226),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_183),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_193),
.C(n_185),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_206),
.B1(n_200),
.B2(n_218),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_265),
.B1(n_239),
.B2(n_229),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_267),
.C(n_268),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_189),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_238),
.C(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_230),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_247),
.B(n_239),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_282),
.B(n_184),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_244),
.B(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_283),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_232),
.B(n_237),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_234),
.C(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_262),
.C(n_267),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_234),
.B1(n_252),
.B2(n_256),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_273),
.B1(n_277),
.B2(n_282),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_296),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_251),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_274),
.B(n_221),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_174),
.C(n_185),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_301),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_295),
.A3(n_289),
.B1(n_290),
.B2(n_296),
.C(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_284),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_174),
.B(n_277),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_304),
.B(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_221),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_180),
.B(n_11),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_279),
.B(n_180),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_293),
.C(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_309),
.B(n_195),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_195),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_313),
.Y(n_315)
);

AO21x2_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_308),
.B(n_192),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_315),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_192),
.B(n_196),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_196),
.Y(n_319)
);


endmodule