module real_jpeg_31402_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_0),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_470),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_1),
.B(n_471),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_47),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_2),
.A2(n_47),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_2),
.A2(n_47),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_108),
.B1(n_183),
.B2(n_188),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_5),
.A2(n_108),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_6),
.Y(n_372)
);

AOI22x1_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_7),
.Y(n_96)
);

OAI22x1_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_96),
.B1(n_154),
.B2(n_158),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_96),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_7),
.B(n_337),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_7),
.A2(n_366),
.A3(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_7),
.B(n_245),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_10),
.A2(n_58),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_10),
.A2(n_58),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_10),
.A2(n_58),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_12),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_259),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_258),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_228),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_19),
.B(n_228),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.C(n_193),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_21),
.B(n_307),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.C(n_101),
.Y(n_21)
);

XOR2x1_ASAP7_75t_L g266 ( 
.A(n_22),
.B(n_63),
.Y(n_266)
);

NAND2x1p5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

NAND2x1p5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_24),
.B(n_54),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_24),
.A2(n_37),
.B(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_24),
.B(n_209),
.Y(n_434)
);

NOR2x1p5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_32),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_36),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_37),
.Y(n_216)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_41),
.Y(n_304)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_45),
.B(n_215),
.Y(n_283)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_53),
.B(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_55),
.Y(n_297)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_90),
.B(n_92),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_64),
.B(n_92),
.Y(n_227)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_64),
.Y(n_248)
);

AO21x2_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_80),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_66),
.Y(n_334)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_71),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_83),
.Y(n_321)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_86),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_87),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_91),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_91),
.Y(n_245)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_92),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_95),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_95),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_96),
.A2(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_96),
.B(n_213),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g330 ( 
.A1(n_96),
.A2(n_331),
.A3(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g349 ( 
.A(n_96),
.B(n_216),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_96),
.B(n_367),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_96),
.B(n_143),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_96),
.B(n_115),
.Y(n_415)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_98),
.Y(n_281)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

XOR2x1_ASAP7_75t_L g265 ( 
.A(n_101),
.B(n_266),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_126),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_102),
.B(n_126),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_113),
.B(n_118),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_103),
.A2(n_205),
.B(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_106),
.Y(n_389)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_107),
.Y(n_388)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_107),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_173),
.B(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_114),
.B(n_121),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_114),
.B(n_176),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_114),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_118),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_118),
.B(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_160),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_127),
.B(n_317),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_153),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_128),
.B(n_318),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_128),
.A2(n_153),
.B(n_161),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_143),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_137),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_146),
.Y(n_380)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_153),
.B(n_233),
.Y(n_232)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_157),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_181),
.B(n_190),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_160),
.B(n_358),
.Y(n_392)
);

NAND2x1p5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_182),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_161),
.B(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_171),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_180),
.B1(n_191),
.B2(n_192),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_172),
.A2(n_191),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_172),
.A2(n_191),
.B1(n_330),
.B2(n_341),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_SL g359 ( 
.A(n_172),
.B(n_330),
.Y(n_359)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_201),
.Y(n_200)
);

BUFx4f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_180),
.B(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_195),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_256),
.C(n_257),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B(n_199),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_197),
.B(n_198),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_197),
.B(n_317),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_199),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

AND2x4_ASAP7_75t_SL g384 ( 
.A(n_200),
.B(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_205),
.B(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_218),
.Y(n_206)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

NAND2x1_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_217),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_212),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_219),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_275),
.Y(n_274)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_224),
.Y(n_293)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_227),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_255),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_250),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_234),
.B(n_249),
.Y(n_230)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_232),
.B(n_358),
.Y(n_357)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_245),
.B(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_245),
.B(n_277),
.Y(n_326)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_247),
.B(n_326),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21x1_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_309),
.B(n_469),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_306),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_262),
.B(n_306),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.C(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_265),
.A2(n_267),
.B1(n_268),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_265),
.Y(n_460)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_271),
.B(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_282),
.C(n_284),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_273),
.B(n_282),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_284),
.B(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_SL g431 ( 
.A(n_285),
.B(n_290),
.Y(n_431)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI31xp33_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_294),
.A3(n_297),
.B(n_298),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_302),
.B(n_305),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_443),
.B(n_463),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_427),
.B(n_441),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_360),
.B(n_426),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_342),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_314),
.B(n_342),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.C(n_328),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_316),
.B(n_325),
.Y(n_424)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_329),
.B(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_356),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_357),
.C(n_359),
.Y(n_440)
);

OAI22x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_347),
.B1(n_354),
.B2(n_355),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_349),
.C(n_350),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_355)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_419),
.B(n_425),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_395),
.B(n_418),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_383),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_383),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_381),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_365),
.B1(n_381),
.B2(n_382),
.Y(n_397)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_373),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_390),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_384),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_391),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_421),
.C(n_422),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_404),
.B(n_417),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_398),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI21x1_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_408),
.B(n_416),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_407),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_420),
.B(n_423),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_440),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_440),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_432),
.C(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_436),
.C(n_438),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_436),
.Y(n_439)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_457),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_451),
.Y(n_465)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_455),
.C(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_454),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_458),
.A2(n_461),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);


endmodule