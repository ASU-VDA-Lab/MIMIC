module fake_jpeg_4348_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_18),
.Y(n_26)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_17),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_19),
.C(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_13),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_8),
.C(n_6),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_27),
.C(n_26),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_6),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_20),
.B1(n_21),
.B2(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_19),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_30),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_35),
.CI(n_36),
.CON(n_39),
.SN(n_39)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_38),
.B1(n_40),
.B2(n_37),
.Y(n_42)
);

BUFx24_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_41),
.B(n_39),
.Y(n_44)
);


endmodule