module fake_jpeg_22889_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_45),
.B1(n_33),
.B2(n_42),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_52),
.B1(n_58),
.B2(n_27),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_45),
.B1(n_33),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_31),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_35),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_33),
.B1(n_20),
.B2(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_65),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_67),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_88),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_20),
.B1(n_27),
.B2(n_23),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_34),
.B(n_29),
.Y(n_119)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_23),
.B1(n_32),
.B2(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_28),
.Y(n_121)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_52),
.B1(n_56),
.B2(n_47),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_99),
.B1(n_106),
.B2(n_107),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_56),
.C(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_13),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_21),
.B(n_22),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_119),
.B(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_47),
.B1(n_42),
.B2(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_22),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_115),
.C(n_39),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_27),
.B1(n_61),
.B2(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_22),
.B1(n_17),
.B2(n_28),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_110),
.B1(n_77),
.B2(n_80),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_17),
.B1(n_28),
.B2(n_31),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_31),
.B1(n_28),
.B2(n_18),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_84),
.C(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_18),
.B1(n_34),
.B2(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_62),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_131),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_126),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_127),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_128),
.A2(n_62),
.B1(n_57),
.B2(n_81),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_139),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_65),
.B(n_30),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_74),
.B(n_83),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_112),
.B(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_138),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_57),
.B1(n_62),
.B2(n_19),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_140),
.B1(n_108),
.B2(n_101),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_39),
.B1(n_36),
.B2(n_41),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_25),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_41),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_148),
.C(n_96),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_36),
.C(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_161),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_149),
.A2(n_97),
.B1(n_99),
.B2(n_98),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_171),
.B1(n_177),
.B2(n_29),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_168),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_106),
.B1(n_107),
.B2(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_95),
.B1(n_103),
.B2(n_94),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_163),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_148),
.C(n_147),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_112),
.B1(n_122),
.B2(n_96),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_176),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_179),
.B(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_5),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_30),
.B(n_36),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_146),
.B(n_10),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_62),
.Y(n_181)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_195),
.B(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_223)
);

BUFx12f_ASAP7_75t_SL g187 ( 
.A(n_169),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_11),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_125),
.C(n_145),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_133),
.C(n_141),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_129),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_197),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_150),
.C(n_137),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_204),
.C(n_160),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_135),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_170),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_29),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_203),
.B1(n_206),
.B2(n_209),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_71),
.B1(n_31),
.B2(n_29),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_0),
.C(n_1),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_178),
.B1(n_173),
.B2(n_161),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_206)
);

INVxp33_ASAP7_75t_SL g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_160),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_2),
.B(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_11),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_175),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_224),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_220),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_171),
.B1(n_168),
.B2(n_162),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_233),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_174),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_232),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_167),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_210),
.C(n_194),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_182),
.B1(n_167),
.B2(n_158),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_182),
.B1(n_172),
.B2(n_155),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_186),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_165),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_252),
.C(n_237),
.Y(n_264)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_190),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_261),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_191),
.C(n_200),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_205),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_257),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_213),
.B(n_206),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_259),
.B(n_163),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_203),
.B(n_209),
.C(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_215),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_232),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_242),
.C(n_247),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_226),
.B1(n_220),
.B2(n_230),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_274),
.B1(n_251),
.B2(n_6),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_278),
.B(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_231),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_223),
.B(n_231),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_275),
.B1(n_251),
.B2(n_12),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_219),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_246),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_204),
.Y(n_273)
);

OAI21x1_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_259),
.B(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_257),
.B1(n_253),
.B2(n_252),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_217),
.B(n_225),
.C(n_180),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_294),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_253),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_264),
.C(n_269),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_259),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_245),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_9),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_266),
.B1(n_273),
.B2(n_13),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_305),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_275),
.B1(n_265),
.B2(n_272),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.C(n_292),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_273),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_306),
.B(n_307),
.Y(n_316)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_304),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_14),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_290),
.C(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_15),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_291),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_285),
.B(n_9),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_308),
.B(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_306),
.B(n_304),
.C(n_293),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_323),
.B1(n_324),
.B2(n_310),
.Y(n_327)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_327),
.C(n_318),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_325),
.B1(n_312),
.B2(n_326),
.Y(n_330)
);

OAI321xp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_314),
.A3(n_15),
.B1(n_8),
.B2(n_7),
.C(n_6),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_6),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_7),
.C(n_8),
.Y(n_333)
);


endmodule