module real_aes_651_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_503;
wire n_792;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_554;
wire n_475;
wire n_798;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g700 ( .A(n_0), .B(n_701), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_1), .Y(n_501) );
AO222x2_ASAP7_75t_SL g572 ( .A1(n_2), .A2(n_33), .B1(n_160), .B2(n_427), .C1(n_443), .C2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_3), .A2(n_24), .B1(n_349), .B2(n_410), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_4), .A2(n_242), .B1(n_451), .B2(n_462), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_5), .A2(n_177), .B1(n_446), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_6), .A2(n_27), .B1(n_499), .B2(n_577), .Y(n_576) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_7), .A2(n_194), .B1(n_310), .B2(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g752 ( .A(n_7), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_8), .A2(n_147), .B1(n_539), .B2(n_565), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_9), .A2(n_137), .B1(n_478), .B2(n_536), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_10), .A2(n_254), .B1(n_632), .B2(n_699), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_11), .A2(n_247), .B1(n_698), .B2(n_699), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_12), .A2(n_268), .B1(n_467), .B2(n_547), .Y(n_558) );
AO22x1_ASAP7_75t_L g765 ( .A1(n_13), .A2(n_201), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_14), .A2(n_78), .B1(n_451), .B2(n_549), .Y(n_675) );
OA22x2_ASAP7_75t_L g676 ( .A1(n_15), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_15), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_16), .A2(n_197), .B1(n_464), .B2(n_465), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_17), .A2(n_30), .B1(n_547), .B2(n_549), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_18), .A2(n_45), .B1(n_365), .B2(n_369), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_19), .A2(n_105), .B1(n_451), .B2(n_462), .Y(n_659) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_20), .A2(n_76), .B1(n_310), .B2(n_311), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_20), .B(n_751), .Y(n_750) );
XOR2x2_ASAP7_75t_L g299 ( .A(n_21), .B(n_300), .Y(n_299) );
XOR2xp5_ASAP7_75t_SL g519 ( .A(n_21), .B(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_22), .A2(n_56), .B1(n_462), .B2(n_547), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_23), .A2(n_161), .B1(n_451), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_25), .A2(n_178), .B1(n_454), .B2(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_26), .A2(n_54), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_28), .A2(n_211), .B1(n_464), .B2(n_465), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_29), .A2(n_74), .B1(n_453), .B2(n_454), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_31), .A2(n_59), .B1(n_338), .B2(n_342), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_32), .A2(n_175), .B1(n_400), .B2(n_402), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_34), .A2(n_71), .B1(n_467), .B2(n_468), .Y(n_685) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_35), .A2(n_239), .B1(n_277), .B2(n_481), .C1(n_482), .C2(n_533), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_36), .A2(n_183), .B1(n_454), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_37), .A2(n_272), .B1(n_303), .B2(n_324), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_38), .A2(n_221), .B1(n_464), .B2(n_465), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_39), .A2(n_95), .B1(n_450), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_40), .A2(n_248), .B1(n_462), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_41), .A2(n_253), .B1(n_402), .B2(n_594), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_42), .A2(n_130), .B1(n_451), .B2(n_462), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_43), .A2(n_174), .B1(n_352), .B2(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_44), .A2(n_192), .B1(n_453), .B2(n_517), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_46), .A2(n_123), .B1(n_481), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_47), .A2(n_48), .B1(n_476), .B2(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_49), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_50), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_51), .A2(n_186), .B1(n_478), .B2(n_536), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_52), .A2(n_60), .B1(n_361), .B2(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_53), .A2(n_267), .B1(n_642), .B2(n_644), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_55), .A2(n_112), .B1(n_405), .B2(n_591), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_57), .B(n_533), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_58), .A2(n_282), .B1(n_530), .B2(n_563), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_61), .A2(n_216), .B1(n_426), .B2(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_62), .A2(n_203), .B1(n_392), .B2(n_394), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_63), .A2(n_172), .B1(n_409), .B2(n_410), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_64), .A2(n_117), .B1(n_424), .B2(n_427), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_65), .A2(n_98), .B1(n_409), .B2(n_577), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_66), .A2(n_219), .B1(n_468), .B2(n_549), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_67), .A2(n_79), .B1(n_371), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_68), .A2(n_145), .B1(n_621), .B2(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_69), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_70), .A2(n_109), .B1(n_377), .B2(n_380), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_72), .A2(n_143), .B1(n_304), .B2(n_468), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_73), .A2(n_90), .B1(n_397), .B2(n_773), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_75), .A2(n_92), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_77), .A2(n_124), .B1(n_539), .B2(n_565), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_80), .A2(n_263), .B1(n_530), .B2(n_531), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_81), .A2(n_280), .B1(n_464), .B2(n_465), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_82), .A2(n_168), .B1(n_365), .B2(n_369), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_83), .A2(n_144), .B1(n_329), .B2(n_333), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_84), .A2(n_115), .B1(n_436), .B2(n_615), .Y(n_614) );
INVx3_ASAP7_75t_L g310 ( .A(n_85), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_86), .A2(n_164), .B1(n_338), .B2(n_436), .Y(n_435) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_87), .A2(n_433), .B1(n_455), .B2(n_456), .Y(n_432) );
INVx1_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_88), .A2(n_135), .B1(n_334), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_89), .A2(n_127), .B1(n_404), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_91), .A2(n_245), .B1(n_358), .B2(n_361), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_93), .A2(n_150), .B1(n_369), .B2(n_448), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_94), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_96), .A2(n_214), .B1(n_338), .B2(n_342), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_97), .A2(n_191), .B1(n_632), .B2(n_633), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_99), .A2(n_180), .B1(n_467), .B2(n_468), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_100), .B(n_422), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_101), .A2(n_114), .B1(n_348), .B2(n_352), .Y(n_347) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_102), .B(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_103), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_104), .A2(n_218), .B1(n_530), .B2(n_531), .Y(n_653) );
INVx1_ASAP7_75t_SL g319 ( .A(n_106), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_106), .B(n_138), .Y(n_753) );
INVx1_ASAP7_75t_L g726 ( .A(n_107), .Y(n_726) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_108), .A2(n_118), .B1(n_241), .B2(n_374), .C1(n_377), .C2(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g292 ( .A(n_110), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_111), .A2(n_281), .B1(n_468), .B2(n_544), .Y(n_543) );
XOR2x2_ASAP7_75t_L g458 ( .A(n_113), .B(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_116), .A2(n_182), .B1(n_402), .B2(n_594), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_119), .A2(n_136), .B1(n_544), .B2(n_547), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_120), .A2(n_134), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_121), .A2(n_224), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_122), .A2(n_285), .B1(n_397), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_125), .A2(n_167), .B1(n_427), .B2(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_126), .A2(n_255), .B1(n_478), .B2(n_536), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_128), .A2(n_229), .B1(n_594), .B2(n_596), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_129), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_131), .A2(n_276), .B1(n_441), .B2(n_473), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_132), .A2(n_237), .B1(n_467), .B2(n_468), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_133), .B(n_414), .Y(n_413) );
AO22x2_ASAP7_75t_L g322 ( .A1(n_138), .A2(n_205), .B1(n_310), .B2(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_139), .A2(n_199), .B1(n_422), .B2(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_140), .B(n_533), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_141), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_142), .B(n_701), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_146), .A2(n_757), .B1(n_781), .B2(n_782), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_146), .Y(n_782) );
XOR2xp5_ASAP7_75t_L g693 ( .A(n_148), .B(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_149), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_151), .B(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_152), .A2(n_264), .B1(n_418), .B2(n_420), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_153), .A2(n_249), .B1(n_304), .B2(n_621), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_154), .A2(n_223), .B1(n_578), .B2(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g320 ( .A(n_155), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_156), .A2(n_262), .B1(n_348), .B2(n_635), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_157), .A2(n_176), .B1(n_325), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_158), .A2(n_278), .B1(n_404), .B2(n_405), .Y(n_403) );
XNOR2xp5_ASAP7_75t_L g488 ( .A(n_159), .B(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_162), .A2(n_244), .B1(n_476), .B2(n_478), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_163), .A2(n_189), .B1(n_464), .B2(n_465), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_165), .B(n_484), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_166), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_169), .A2(n_271), .B1(n_352), .B2(n_409), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_170), .A2(n_230), .B1(n_326), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_171), .A2(n_193), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_173), .A2(n_206), .B1(n_464), .B2(n_465), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_179), .Y(n_722) );
XNOR2x1_ASAP7_75t_L g664 ( .A(n_181), .B(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_184), .A2(n_208), .B1(n_470), .B2(n_621), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_185), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_187), .A2(n_220), .B1(n_536), .B2(n_537), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_188), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_190), .A2(n_265), .B1(n_536), .B2(n_537), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_195), .A2(n_257), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_196), .A2(n_243), .B1(n_349), .B2(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_198), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g550 ( .A(n_200), .Y(n_550) );
INVx1_ASAP7_75t_L g801 ( .A(n_202), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_204), .A2(n_246), .B1(n_358), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_207), .A2(n_256), .B1(n_530), .B2(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_209), .B(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_210), .A2(n_251), .B1(n_333), .B2(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_212), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_213), .B(n_374), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_215), .Y(n_714) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_217), .A2(n_570), .B(n_597), .Y(n_569) );
INVx1_ASAP7_75t_L g599 ( .A(n_217), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_222), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_225), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g748 ( .A(n_225), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_226), .A2(n_258), .B1(n_481), .B2(n_482), .Y(n_480) );
AO22x2_ASAP7_75t_L g553 ( .A1(n_227), .A2(n_554), .B1(n_567), .B2(n_568), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_227), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_228), .A2(n_269), .B1(n_381), .B2(n_441), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_231), .A2(n_240), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g289 ( .A(n_232), .Y(n_289) );
AND2x2_ASAP7_75t_R g784 ( .A(n_232), .B(n_748), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_233), .A2(n_236), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_234), .A2(n_283), .B1(n_450), .B2(n_621), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_235), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_238), .A2(n_624), .B1(n_625), .B2(n_645), .Y(n_623) );
INVx1_ASAP7_75t_L g645 ( .A(n_238), .Y(n_645) );
INVxp67_ASAP7_75t_L g294 ( .A(n_250), .Y(n_294) );
XNOR2x1_ASAP7_75t_L g607 ( .A(n_252), .B(n_608), .Y(n_607) );
XOR2xp5_ASAP7_75t_L g661 ( .A(n_252), .B(n_608), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_259), .B(n_484), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_260), .A2(n_270), .B1(n_451), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_261), .A2(n_273), .B1(n_349), .B2(n_731), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_266), .A2(n_287), .B1(n_295), .B2(n_754), .C(n_755), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_274), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_275), .A2(n_279), .B1(n_482), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_284), .Y(n_709) );
NOR2x1_ASAP7_75t_R g287 ( .A(n_288), .B(n_290), .Y(n_287) );
OR2x2_ASAP7_75t_L g805 ( .A(n_288), .B(n_291), .Y(n_805) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_289), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI21xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_601), .B(n_745), .Y(n_295) );
OR2x2_ASAP7_75t_L g754 ( .A(n_296), .B(n_601), .Y(n_754) );
AOI22xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_522), .B1(n_523), .B2(n_600), .Y(n_296) );
INVx1_ASAP7_75t_L g600 ( .A(n_297), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_385), .B1(n_519), .B2(n_521), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_300), .Y(n_520) );
NAND4xp75_ASAP7_75t_SL g300 ( .A(n_301), .B(n_336), .C(n_356), .D(n_373), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_328), .Y(n_301) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx3_ASAP7_75t_SL g404 ( .A(n_305), .Y(n_404) );
INVx2_ASAP7_75t_L g446 ( .A(n_305), .Y(n_446) );
INVx3_ASAP7_75t_L g470 ( .A(n_305), .Y(n_470) );
INVx2_ASAP7_75t_SL g513 ( .A(n_305), .Y(n_513) );
INVx2_ASAP7_75t_SL g741 ( .A(n_305), .Y(n_741) );
INVx8_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_315), .Y(n_306) );
AND2x4_ASAP7_75t_L g331 ( .A(n_307), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_307), .B(n_351), .Y(n_360) );
AND2x2_ASAP7_75t_L g376 ( .A(n_307), .B(n_344), .Y(n_376) );
AND2x6_ASAP7_75t_L g462 ( .A(n_307), .B(n_351), .Y(n_462) );
AND2x2_ASAP7_75t_L g467 ( .A(n_307), .B(n_332), .Y(n_467) );
AND2x4_ASAP7_75t_L g533 ( .A(n_307), .B(n_344), .Y(n_533) );
AND2x2_ASAP7_75t_L g544 ( .A(n_307), .B(n_332), .Y(n_544) );
AND2x2_ASAP7_75t_L g549 ( .A(n_307), .B(n_315), .Y(n_549) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g327 ( .A(n_309), .B(n_312), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
INVx2_ASAP7_75t_L g311 ( .A(n_310), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_310), .Y(n_314) );
OAI22x1_ASAP7_75t_L g317 ( .A1(n_310), .A2(n_318), .B1(n_319), .B2(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_310), .Y(n_318) );
INVx1_ASAP7_75t_L g323 ( .A(n_310), .Y(n_323) );
INVxp67_ASAP7_75t_L g355 ( .A(n_312), .Y(n_355) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g340 ( .A(n_313), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g326 ( .A(n_315), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g334 ( .A(n_315), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g363 ( .A(n_315), .B(n_340), .Y(n_363) );
AND2x6_ASAP7_75t_L g451 ( .A(n_315), .B(n_340), .Y(n_451) );
AND2x4_ASAP7_75t_L g468 ( .A(n_315), .B(n_335), .Y(n_468) );
AND2x2_ASAP7_75t_L g547 ( .A(n_315), .B(n_327), .Y(n_547) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x2_ASAP7_75t_L g351 ( .A(n_316), .B(n_322), .Y(n_351) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g332 ( .A(n_317), .B(n_321), .Y(n_332) );
AND2x2_ASAP7_75t_L g344 ( .A(n_317), .B(n_322), .Y(n_344) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g724 ( .A(n_325), .Y(n_724) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_326), .Y(n_517) );
BUFx3_ASAP7_75t_L g585 ( .A(n_326), .Y(n_585) );
AND2x4_ASAP7_75t_L g350 ( .A(n_327), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g379 ( .A(n_327), .B(n_332), .Y(n_379) );
AND2x2_ASAP7_75t_L g481 ( .A(n_327), .B(n_351), .Y(n_481) );
AND2x4_ASAP7_75t_L g530 ( .A(n_327), .B(n_332), .Y(n_530) );
AND2x2_ASAP7_75t_L g565 ( .A(n_327), .B(n_351), .Y(n_565) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g396 ( .A(n_330), .Y(n_396) );
INVx2_ASAP7_75t_L g509 ( .A(n_330), .Y(n_509) );
INVx2_ASAP7_75t_L g638 ( .A(n_330), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_330), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
INVx3_ASAP7_75t_L g773 ( .A(n_330), .Y(n_773) );
INVx6_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g453 ( .A(n_331), .Y(n_453) );
BUFx3_ASAP7_75t_L g588 ( .A(n_331), .Y(n_588) );
AND2x2_ASAP7_75t_L g339 ( .A(n_332), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g536 ( .A(n_332), .B(n_340), .Y(n_536) );
BUFx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g398 ( .A(n_334), .Y(n_398) );
BUFx3_ASAP7_75t_L g454 ( .A(n_334), .Y(n_454) );
AND2x4_ASAP7_75t_L g371 ( .A(n_335), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g465 ( .A(n_335), .B(n_372), .Y(n_465) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_335), .B(n_384), .Y(n_531) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_335), .B(n_384), .Y(n_563) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_347), .Y(n_336) );
BUFx6f_ASAP7_75t_SL g409 ( .A(n_338), .Y(n_409) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g477 ( .A(n_339), .Y(n_477) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_339), .Y(n_615) );
AND2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_351), .Y(n_368) );
AND2x2_ASAP7_75t_L g464 ( .A(n_340), .B(n_351), .Y(n_464) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_341), .Y(n_346) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g412 ( .A(n_343), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_343), .Y(n_437) );
BUFx6f_ASAP7_75t_SL g578 ( .A(n_343), .Y(n_578) );
BUFx3_ASAP7_75t_L g780 ( .A(n_343), .Y(n_780) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x4_ASAP7_75t_L g354 ( .A(n_344), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g478 ( .A(n_344), .B(n_345), .Y(n_478) );
AND2x2_ASAP7_75t_L g482 ( .A(n_344), .B(n_355), .Y(n_482) );
AND2x2_ASAP7_75t_L g537 ( .A(n_344), .B(n_345), .Y(n_537) );
AND2x2_ASAP7_75t_L g539 ( .A(n_344), .B(n_355), .Y(n_539) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g504 ( .A(n_348), .Y(n_504) );
BUFx4f_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g573 ( .A(n_349), .Y(n_573) );
BUFx2_ASAP7_75t_L g762 ( .A(n_349), .Y(n_762) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g426 ( .A(n_350), .Y(n_426) );
BUFx2_ASAP7_75t_L g613 ( .A(n_350), .Y(n_613) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
INVx2_ASAP7_75t_L g439 ( .A(n_353), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_353), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
INVx2_ASAP7_75t_SL g635 ( .A(n_353), .Y(n_635) );
INVx1_ASAP7_75t_L g731 ( .A(n_353), .Y(n_731) );
INVx6_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_364), .Y(n_356) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g591 ( .A(n_359), .Y(n_591) );
INVx2_ASAP7_75t_L g643 ( .A(n_359), .Y(n_643) );
INVx2_ASAP7_75t_L g737 ( .A(n_359), .Y(n_737) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g393 ( .A(n_360), .Y(n_393) );
BUFx2_ASAP7_75t_L g450 ( .A(n_360), .Y(n_450) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g394 ( .A(n_362), .Y(n_394) );
INVx2_ASAP7_75t_SL g592 ( .A(n_362), .Y(n_592) );
INVx2_ASAP7_75t_L g621 ( .A(n_362), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_362), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx2_ASAP7_75t_L g771 ( .A(n_362), .Y(n_771) );
INVx8_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g719 ( .A(n_366), .Y(n_719) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_366), .Y(n_766) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g595 ( .A(n_367), .Y(n_595) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_368), .Y(n_448) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
INVx2_ASAP7_75t_L g596 ( .A(n_370), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_370), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_716) );
INVx5_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g767 ( .A(n_371), .Y(n_767) );
BUFx2_ASAP7_75t_L g799 ( .A(n_374), .Y(n_799) );
INVx4_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_SL g416 ( .A(n_375), .Y(n_416) );
INVx3_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
INVx4_ASAP7_75t_SL g484 ( .A(n_375), .Y(n_484) );
INVx3_ASAP7_75t_L g629 ( .A(n_375), .Y(n_629) );
BUFx2_ASAP7_75t_L g702 ( .A(n_375), .Y(n_702) );
INVx6_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g494 ( .A(n_378), .Y(n_494) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
BUFx3_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g473 ( .A(n_382), .Y(n_473) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx12f_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
INVx1_ASAP7_75t_SL g521 ( .A(n_385), .Y(n_521) );
XNOR2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_485), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_429), .B2(n_430), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
XOR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_428), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_407), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .C(n_399), .D(n_403), .Y(n_390) );
INVx1_ASAP7_75t_L g713 ( .A(n_392), .Y(n_713) );
BUFx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g710 ( .A(n_397), .Y(n_710) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g775 ( .A(n_406), .Y(n_775) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_413), .C(n_417), .D(n_423), .Y(n_407) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_411), .A2(n_497), .B1(n_498), .B2(n_501), .Y(n_496) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_415), .A2(n_492), .B1(n_493), .B2(n_494), .C(n_495), .Y(n_491) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
INVx1_ASAP7_75t_L g698 ( .A(n_419), .Y(n_698) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g699 ( .A(n_422), .Y(n_699) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OA22x2_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_457), .B2(n_458), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g456 ( .A(n_433), .Y(n_456) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_444), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .C(n_440), .D(n_442), .Y(n_434) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_441), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .C(n_449), .D(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g581 ( .A(n_446), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_457), .A2(n_458), .B1(n_488), .B2(n_518), .Y(n_487) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_479), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .C(n_466), .D(n_469), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
BUFx2_ASAP7_75t_L g633 ( .A(n_473), .Y(n_633) );
INVx4_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g500 ( .A(n_477), .Y(n_500) );
INVx2_ASAP7_75t_L g734 ( .A(n_477), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g518 ( .A(n_488), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_506), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_496), .C(n_502), .Y(n_490) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_517), .Y(n_644) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
XNOR2xp5_ASAP7_75t_SL g523 ( .A(n_524), .B(n_551), .Y(n_523) );
INVx3_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
XOR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_550), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_540), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_532), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_569), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g568 ( .A(n_554), .Y(n_568) );
NOR2xp67_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .C(n_558), .D(n_559), .Y(n_555) );
NAND4xp25_ASAP7_75t_SL g560 ( .A(n_561), .B(n_562), .C(n_564), .D(n_566), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_579), .C(n_589), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
NOR4xp25_ASAP7_75t_L g597 ( .A(n_572), .B(n_574), .C(n_580), .D(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
BUFx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B1(n_583), .B2(n_586), .C(n_587), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_581), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_589), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_691), .B1(n_743), .B2(n_744), .Y(n_601) );
INVx1_ASAP7_75t_L g744 ( .A(n_602), .Y(n_744) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_663), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_622), .B2(n_662), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_607), .A2(n_648), .B1(n_649), .B2(n_661), .Y(n_647) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_616), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .C(n_612), .D(n_614), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .C(n_619), .D(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_646), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_636), .Y(n_625) );
NAND4xp25_ASAP7_75t_SL g626 ( .A(n_627), .B(n_630), .C(n_631), .D(n_634), .Y(n_626) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .C(n_640), .D(n_641), .Y(n_636) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
NAND4xp25_ASAP7_75t_SL g651 ( .A(n_652), .B(n_653), .C(n_654), .D(n_655), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .C(n_659), .D(n_660), .Y(n_656) );
AO22x2_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_676), .B1(n_689), .B2(n_690), .Y(n_663) );
INVx1_ASAP7_75t_L g689 ( .A(n_664), .Y(n_689) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_671), .Y(n_665) );
NAND4xp25_ASAP7_75t_SL g666 ( .A(n_667), .B(n_668), .C(n_669), .D(n_670), .Y(n_666) );
NAND4xp25_ASAP7_75t_SL g671 ( .A(n_672), .B(n_673), .C(n_674), .D(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g690 ( .A(n_676), .Y(n_690) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .C(n_683), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .C(n_687), .D(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g743 ( .A(n_691), .Y(n_743) );
OAI22xp33_ASAP7_75t_R g691 ( .A1(n_692), .A2(n_693), .B1(n_725), .B2(n_742), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .C(n_715), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_703), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_700), .Y(n_696) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_711), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_721), .Y(n_715) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g742 ( .A(n_725), .Y(n_742) );
XNOR2x2_ASAP7_75t_SL g725 ( .A(n_726), .B(n_727), .Y(n_725) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_735), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_732), .D(n_733), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .C(n_739), .D(n_740), .Y(n_735) );
INVx4_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_747), .B(n_750), .Y(n_804) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
OAI222xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_783), .B1(n_785), .B2(n_801), .C1(n_802), .C2(n_805), .Y(n_755) );
INVx1_ASAP7_75t_L g781 ( .A(n_757), .Y(n_781) );
NAND5xp2_ASAP7_75t_L g757 ( .A(n_758), .B(n_763), .C(n_764), .D(n_768), .E(n_776), .Y(n_757) );
INVxp33_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .C(n_774), .Y(n_769) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_775), .Y(n_792) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx6f_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
XNOR2x1_ASAP7_75t_L g787 ( .A(n_788), .B(n_801), .Y(n_787) );
NOR2xp67_ASAP7_75t_L g788 ( .A(n_789), .B(n_795), .Y(n_788) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .C(n_793), .D(n_794), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_798), .D(n_800), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
CKINVDCx6p67_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
endmodule