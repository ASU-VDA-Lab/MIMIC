module fake_jpeg_2069_n_522 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_522);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_522;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_29),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_66),
.B(n_97),
.Y(n_113)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_80),
.Y(n_141)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_1),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_98),
.B(n_44),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_115),
.B(n_137),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_34),
.B1(n_47),
.B2(n_43),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_117),
.A2(n_153),
.B1(n_32),
.B2(n_43),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_47),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_123),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_55),
.A2(n_33),
.B1(n_48),
.B2(n_47),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_128),
.A2(n_150),
.B1(n_159),
.B2(n_61),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_83),
.B(n_36),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_71),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_32),
.B1(n_91),
.B2(n_86),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_52),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_60),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_89),
.A2(n_33),
.B1(n_48),
.B2(n_28),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_57),
.A2(n_33),
.B1(n_48),
.B2(n_44),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_58),
.B1(n_99),
.B2(n_95),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_161),
.A2(n_143),
.B1(n_138),
.B2(n_126),
.Y(n_261)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_36),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_172),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_167),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g254 ( 
.A(n_171),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_50),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_176),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_199),
.B1(n_203),
.B2(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_180),
.Y(n_227)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_75),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_198),
.B1(n_68),
.B2(n_84),
.Y(n_224)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_111),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_189),
.Y(n_229)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_50),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_125),
.B(n_35),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_101),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_196),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_118),
.A2(n_102),
.B1(n_54),
.B2(n_69),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_201),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_110),
.Y(n_201)
);

CKINVDCx6p67_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_204),
.Y(n_231)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_239)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

BUFx16f_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_101),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_35),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_119),
.Y(n_246)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_138),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_165),
.A2(n_128),
.B1(n_150),
.B2(n_159),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_218),
.A2(n_40),
.B1(n_51),
.B2(n_45),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_82),
.C(n_156),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_233),
.C(n_252),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_224),
.A2(n_228),
.B1(n_251),
.B2(n_51),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_157),
.B1(n_142),
.B2(n_134),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_226),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_22),
.B1(n_25),
.B2(n_39),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_80),
.B(n_25),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_233),
.A2(n_241),
.B(n_199),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_80),
.B(n_22),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_155),
.B1(n_158),
.B2(n_146),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_253),
.B1(n_263),
.B2(n_185),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_142),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_252),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_176),
.A2(n_96),
.B1(n_88),
.B2(n_134),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_136),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_168),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_174),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_164),
.Y(n_277)
);

AO21x2_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_45),
.B(n_59),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_200),
.A2(n_87),
.B1(n_94),
.B2(n_85),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_175),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_265),
.B(n_298),
.Y(n_334)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

BUFx2_ASAP7_75t_SL g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_162),
.A3(n_171),
.B1(n_192),
.B2(n_208),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_270),
.B(n_307),
.C(n_263),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_136),
.B1(n_143),
.B2(n_183),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_271),
.A2(n_278),
.B1(n_286),
.B2(n_292),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_280),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_296),
.C(n_235),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_224),
.A2(n_202),
.B(n_193),
.C(n_206),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_276),
.A2(n_232),
.B(n_254),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_287),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_93),
.B1(n_100),
.B2(n_81),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_231),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_282),
.B(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_207),
.B(n_184),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_284),
.A2(n_293),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_220),
.A2(n_196),
.B1(n_46),
.B2(n_49),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_49),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_242),
.A2(n_39),
.B1(n_46),
.B2(n_209),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_288),
.A2(n_297),
.B1(n_239),
.B2(n_217),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_225),
.B(n_202),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_255),
.C(n_240),
.Y(n_341)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_220),
.B(n_197),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_301),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_231),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_223),
.B(n_59),
.C(n_98),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_236),
.A2(n_45),
.B1(n_51),
.B2(n_40),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_1),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_238),
.B(n_1),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_299),
.B(n_300),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_1),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_2),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_2),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_3),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_3),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_SL g307 ( 
.A(n_241),
.B(n_3),
.C(n_5),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_226),
.B(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_245),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_313),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_277),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_315),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_341),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_269),
.A2(n_226),
.B1(n_262),
.B2(n_253),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_346),
.B1(n_271),
.B2(n_284),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_279),
.A2(n_244),
.B1(n_245),
.B2(n_262),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_324),
.A2(n_332),
.B1(n_335),
.B2(n_342),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_329),
.Y(n_361)
);

NOR2x1p5_ASAP7_75t_SL g329 ( 
.A(n_266),
.B(n_244),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_286),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_254),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_284),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_279),
.A2(n_262),
.B1(n_222),
.B2(n_257),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_333),
.A2(n_343),
.B(n_344),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_279),
.A2(n_222),
.B1(n_257),
.B2(n_255),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_296),
.C(n_274),
.Y(n_358)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_272),
.A2(n_237),
.B1(n_230),
.B2(n_240),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_293),
.A2(n_237),
.B(n_250),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_282),
.A2(n_250),
.B(n_230),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_274),
.A2(n_249),
.B1(n_248),
.B2(n_235),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_295),
.B(n_276),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_355),
.B1(n_357),
.B2(n_372),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_341),
.B(n_289),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_358),
.C(n_375),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_308),
.B1(n_306),
.B2(n_291),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_275),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_364),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_362),
.C(n_369),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_273),
.C(n_280),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_317),
.A2(n_315),
.B1(n_314),
.B2(n_310),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_346),
.B1(n_331),
.B2(n_344),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_302),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_301),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_379),
.Y(n_405)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_311),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_373),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_278),
.C(n_249),
.Y(n_369)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_328),
.A2(n_295),
.B(n_304),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_371),
.A2(n_335),
.B(n_342),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_318),
.A2(n_292),
.B1(n_281),
.B2(n_288),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_327),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_292),
.B1(n_307),
.B2(n_297),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_380),
.B1(n_312),
.B2(n_337),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_248),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_348),
.C(n_320),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_292),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_318),
.A2(n_292),
.B1(n_268),
.B2(n_254),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_347),
.B(n_5),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_381),
.B(n_326),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_328),
.A2(n_264),
.B(n_6),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_368),
.A2(n_325),
.B1(n_333),
.B2(n_324),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_396),
.B1(n_399),
.B2(n_402),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_363),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_390),
.Y(n_427)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_362),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_376),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_391),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_395),
.Y(n_433)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_326),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_370),
.A2(n_352),
.B1(n_349),
.B2(n_361),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_397),
.B(n_350),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_398),
.A2(n_371),
.B(n_380),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_361),
.A2(n_316),
.B1(n_332),
.B2(n_329),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_329),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_337),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_374),
.A2(n_340),
.B1(n_339),
.B2(n_338),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_334),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_406),
.Y(n_435)
);

AOI22x1_ASAP7_75t_L g407 ( 
.A1(n_354),
.A2(n_313),
.B1(n_320),
.B2(n_338),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_264),
.B1(n_8),
.B2(n_9),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_382),
.Y(n_409)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_312),
.C(n_322),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_378),
.C(n_365),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_359),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_401),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_417),
.C(n_418),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_373),
.C(n_369),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_350),
.C(n_377),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_421),
.B(n_429),
.Y(n_445)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_423),
.B(n_436),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_426),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_379),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_428),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_412),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_351),
.C(n_360),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_437),
.C(n_405),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_385),
.A2(n_366),
.B(n_359),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_434),
.Y(n_452)
);

BUFx24_ASAP7_75t_SL g432 ( 
.A(n_395),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_432),
.Y(n_442)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_264),
.C(n_8),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_389),
.B1(n_411),
.B2(n_404),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_439),
.A2(n_441),
.B1(n_443),
.B2(n_447),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_388),
.B1(n_407),
.B2(n_435),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_425),
.A2(n_420),
.B1(n_419),
.B2(n_396),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_425),
.A2(n_403),
.B1(n_385),
.B2(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_410),
.C(n_392),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_457),
.C(n_459),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_420),
.A2(n_403),
.B1(n_405),
.B2(n_400),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_427),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_418),
.C(n_430),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_402),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_458),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_399),
.C(n_383),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_461),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_414),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_443),
.A2(n_419),
.B1(n_415),
.B2(n_424),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_463),
.A2(n_464),
.B1(n_452),
.B2(n_453),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_447),
.A2(n_423),
.B1(n_436),
.B2(n_426),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_442),
.B(n_416),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_466),
.B(n_472),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_437),
.C(n_438),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_471),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_5),
.C(n_9),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_9),
.C(n_10),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_10),
.C(n_11),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_10),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_445),
.B1(n_458),
.B2(n_450),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_476),
.A2(n_449),
.B1(n_13),
.B2(n_14),
.Y(n_501)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_479),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_446),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_484),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_459),
.C(n_446),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_482),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_442),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_453),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_486),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_451),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_487),
.B(n_490),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_471),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_489),
.A2(n_474),
.B1(n_472),
.B2(n_475),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_481),
.C(n_486),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_488),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_476),
.A2(n_454),
.B(n_473),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_497),
.B(n_499),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_454),
.B(n_483),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_448),
.B(n_444),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_501),
.B(n_449),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_506),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_485),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_509),
.B(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_10),
.C(n_13),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_15),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_15),
.B(n_16),
.Y(n_509)
);

AOI31xp33_ASAP7_75t_L g514 ( 
.A1(n_510),
.A2(n_511),
.A3(n_513),
.B(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_496),
.Y(n_511)
);

OAI21x1_ASAP7_75t_SL g518 ( 
.A1(n_514),
.A2(n_516),
.B(n_502),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_512),
.A2(n_503),
.B(n_494),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_515),
.B(n_499),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_512),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_517),
.A2(n_518),
.B(n_505),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_495),
.C(n_501),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_495),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_17),
.B(n_15),
.Y(n_522)
);


endmodule