module fake_jpeg_25684_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_3),
.B(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_39),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_46),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_59),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_43),
.B1(n_44),
.B2(n_26),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_27),
.B1(n_21),
.B2(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_70),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_35),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_26),
.B1(n_28),
.B2(n_25),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_86),
.B1(n_90),
.B2(n_96),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_20),
.B1(n_24),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_71),
.B1(n_61),
.B2(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_108),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_45),
.B1(n_27),
.B2(n_21),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_80),
.B1(n_53),
.B2(n_61),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_59),
.B(n_57),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_88),
.CON(n_155),
.SN(n_155)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_133),
.B1(n_134),
.B2(n_92),
.Y(n_154)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_135),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_45),
.B1(n_52),
.B2(n_21),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_45),
.B(n_57),
.C(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_77),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_77),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_105),
.B1(n_96),
.B2(n_104),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_145),
.B(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_96),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_149),
.B1(n_153),
.B2(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_83),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_96),
.B1(n_101),
.B2(n_108),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_83),
.C(n_89),
.Y(n_150)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_14),
.C(n_5),
.D(n_6),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_98),
.B1(n_93),
.B2(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_132),
.B1(n_116),
.B2(n_120),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_110),
.B1(n_109),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_156),
.A2(n_120),
.B1(n_127),
.B2(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_106),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_111),
.B1(n_3),
.B2(n_4),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_2),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_164),
.B1(n_177),
.B2(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_127),
.C(n_122),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_173),
.C(n_140),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_14),
.C(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_131),
.C(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_121),
.B1(n_113),
.B2(n_7),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_113),
.B1(n_6),
.B2(n_8),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_145),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_150),
.B(n_155),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_189),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_139),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_139),
.C(n_141),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_195),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_191),
.B(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_138),
.C(n_145),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_146),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_154),
.C(n_152),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_182),
.B1(n_171),
.B2(n_173),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_163),
.B1(n_168),
.B2(n_188),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_187),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_162),
.B(n_191),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

AO221x1_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_166),
.B1(n_172),
.B2(n_176),
.C(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_202),
.C(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_168),
.B1(n_198),
.B2(n_184),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_2),
.B(n_9),
.C(n_10),
.Y(n_219)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_9),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_210),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_218),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_224),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_212),
.C(n_207),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_219),
.B(n_222),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_213),
.C(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_10),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_204),
.B1(n_206),
.B2(n_212),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_227),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_219),
.B1(n_205),
.B2(n_12),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_240),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_11),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_233),
.B(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_241),
.C(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_245),
.Y(n_247)
);


endmodule