module fake_aes_12009_n_614 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_614);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_614;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g73 ( .A(n_48), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_31), .Y(n_74) );
INVxp67_ASAP7_75t_L g75 ( .A(n_53), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_25), .Y(n_76) );
CKINVDCx14_ASAP7_75t_R g77 ( .A(n_41), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_63), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_11), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_44), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_47), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_51), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_30), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_4), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_8), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_32), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_34), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_6), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_6), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
INVx1_ASAP7_75t_SL g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_59), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_35), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_0), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_22), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_71), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_57), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_5), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_28), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_27), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
NOR2xp67_ASAP7_75t_L g108 ( .A(n_49), .B(n_10), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_64), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_29), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_5), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_70), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_43), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_67), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_82), .B(n_79), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_96), .B(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_74), .A2(n_33), .B(n_69), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_100), .B(n_1), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_100), .B(n_2), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_111), .B(n_3), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_79), .B(n_3), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g137 ( .A(n_103), .B(n_72), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_116), .B(n_4), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_81), .B(n_36), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_80), .B(n_7), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_97), .B(n_7), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_105), .Y(n_149) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_107), .A2(n_37), .B(n_62), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_107), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_80), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_110), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_104), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_131), .A2(n_117), .B1(n_115), .B2(n_86), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_139), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_131), .B(n_112), .C(n_115), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_118), .B(n_109), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_130), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_128), .A2(n_117), .B1(n_86), .B2(n_91), .Y(n_164) );
INVxp33_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_152), .B(n_77), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_118), .B(n_75), .Y(n_170) );
INVxp67_ASAP7_75t_SL g171 ( .A(n_152), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
CKINVDCx11_ASAP7_75t_R g173 ( .A(n_126), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_128), .A2(n_98), .B1(n_91), .B2(n_93), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_120), .B(n_73), .Y(n_175) );
AND2x6_ASAP7_75t_L g176 ( .A(n_124), .B(n_114), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_124), .B(n_99), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_138), .B(n_98), .C(n_93), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_138), .B(n_99), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_120), .B(n_102), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_138), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_124), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_132), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_132), .B(n_95), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_123), .A2(n_113), .B1(n_106), .B2(n_78), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_130), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_137), .B(n_108), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_123), .B(n_101), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_130), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_142), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_129), .B(n_83), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_133), .B(n_92), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_156), .A2(n_9), .B1(n_12), .B2(n_13), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_140), .B(n_65), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_156), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
INVx5_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_133), .B(n_12), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_177), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_136), .B1(n_144), .B2(n_141), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_189), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_171), .B(n_141), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
INVx5_ASAP7_75t_L g218 ( .A(n_207), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_187), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_177), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_177), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_204), .B(n_149), .Y(n_223) );
OR2x6_ASAP7_75t_L g224 ( .A(n_206), .B(n_144), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_160), .B(n_134), .Y(n_225) );
INVxp67_ASAP7_75t_SL g226 ( .A(n_166), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_203), .B(n_134), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_165), .B(n_145), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_177), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_179), .B(n_145), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_179), .B(n_178), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_189), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_177), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_169), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_165), .B(n_148), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_176), .A2(n_149), .B1(n_148), .B2(n_140), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_203), .B(n_146), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_166), .B(n_137), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_169), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_169), .Y(n_246) );
BUFx12f_ASAP7_75t_L g247 ( .A(n_173), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_161), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_176), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_176), .A2(n_143), .B1(n_146), .B2(n_147), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_161), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_202), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_164), .B(n_146), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_158), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_176), .A2(n_146), .B1(n_143), .B2(n_119), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_175), .B(n_143), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_186), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_182), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_176), .B(n_136), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_195), .A2(n_173), .B1(n_208), .B2(n_168), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_186), .B(n_143), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_195), .A2(n_122), .B1(n_154), .B2(n_153), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_157), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_162), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_167), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_190), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_239), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_245), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_230), .B(n_181), .Y(n_274) );
CKINVDCx8_ASAP7_75t_R g275 ( .A(n_261), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_239), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_244), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_265), .A2(n_208), .B1(n_205), .B2(n_159), .C(n_174), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_245), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_231), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_224), .A2(n_190), .B1(n_192), .B2(n_170), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_247), .A2(n_190), .B1(n_207), .B2(n_196), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_230), .B(n_135), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_225), .A2(n_188), .B(n_201), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_244), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_246), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_247), .B(n_188), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_230), .B(n_190), .Y(n_291) );
NAND2xp33_ASAP7_75t_L g292 ( .A(n_218), .B(n_172), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_213), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_234), .B(n_207), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_216), .B(n_190), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_262), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_213), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_212), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_216), .B(n_135), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_234), .B(n_207), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_226), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_224), .A2(n_190), .B1(n_207), .B2(n_211), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_261), .A2(n_188), .B1(n_201), .B2(n_122), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_234), .B(n_158), .Y(n_305) );
NAND2x1_ASAP7_75t_SL g306 ( .A(n_262), .B(n_122), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_224), .A2(n_125), .B1(n_127), .B2(n_135), .C(n_153), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_257), .A2(n_210), .B(n_197), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_234), .B(n_207), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_249), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_228), .A2(n_154), .B(n_127), .C(n_153), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_220), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_220), .B(n_210), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_214), .B(n_154), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_224), .B1(n_261), .B2(n_254), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_276), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_286), .A2(n_243), .B(n_227), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_275), .A2(n_261), .B1(n_264), .B2(n_250), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_275), .A2(n_256), .B1(n_224), .B2(n_241), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_299), .B(n_283), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_254), .B1(n_240), .B2(n_242), .C(n_223), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_276), .Y(n_323) );
CKINVDCx6p67_ASAP7_75t_R g324 ( .A(n_290), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_280), .A2(n_268), .B1(n_267), .B2(n_266), .C(n_258), .Y(n_325) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_287), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_279), .Y(n_327) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_294), .B(n_269), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_296), .A2(n_218), .B1(n_269), .B2(n_221), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_299), .B(n_268), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_302), .A2(n_267), .B1(n_266), .B2(n_218), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_277), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_296), .A2(n_258), .B1(n_259), .B2(n_219), .C(n_233), .Y(n_333) );
OAI211xp5_ASAP7_75t_L g334 ( .A1(n_281), .A2(n_263), .B(n_127), .C(n_125), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_290), .B(n_238), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_283), .B(n_263), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_290), .B(n_221), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_237), .B(n_219), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_277), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_322), .A2(n_307), .B1(n_284), .B2(n_301), .C(n_314), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_319), .A2(n_300), .B1(n_294), .B2(n_309), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_320), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_320), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_315), .A2(n_311), .B1(n_295), .B2(n_294), .C(n_309), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_321), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_317), .A2(n_285), .B(n_298), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_328), .A2(n_309), .B1(n_300), .B2(n_326), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_321), .B(n_300), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_335), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_333), .A2(n_300), .B1(n_309), .B2(n_290), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_330), .B(n_306), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_324), .A2(n_282), .B1(n_291), .B2(n_310), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_290), .B1(n_218), .B2(n_288), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_325), .A2(n_306), .B1(n_305), .B2(n_304), .C(n_125), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_330), .B(n_271), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_336), .A2(n_236), .B1(n_233), .B2(n_232), .C(n_271), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_338), .B(n_288), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_336), .A2(n_232), .B1(n_236), .B2(n_289), .C(n_155), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_334), .A2(n_142), .B(n_155), .C(n_151), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_342), .B(n_289), .Y(n_366) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_332), .B(n_338), .C(n_341), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_345), .B(n_328), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_347), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_349), .B(n_323), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_361), .B(n_342), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_350), .A2(n_340), .B(n_331), .Y(n_372) );
AOI33xp33_ASAP7_75t_L g373 ( .A1(n_346), .A2(n_332), .A3(n_163), .B1(n_329), .B2(n_17), .B3(n_14), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_347), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_345), .A2(n_328), .B1(n_318), .B2(n_335), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_346), .B(n_327), .Y(n_377) );
OAI33xp33_ASAP7_75t_L g378 ( .A1(n_356), .A2(n_163), .A3(n_200), .B1(n_198), .B2(n_185), .B3(n_183), .Y(n_378) );
OAI211xp5_ASAP7_75t_L g379 ( .A1(n_355), .A2(n_155), .B(n_151), .C(n_142), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_339), .B1(n_335), .B2(n_326), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_366), .B(n_121), .Y(n_381) );
OA21x2_ASAP7_75t_L g382 ( .A1(n_367), .A2(n_150), .B(n_121), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_354), .B(n_335), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_353), .B(n_327), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_366), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_353), .B(n_335), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_360), .B(n_339), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_354), .B(n_339), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_352), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_343), .B(n_142), .C(n_151), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_344), .B(n_348), .C(n_363), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_362), .B(n_121), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_358), .A2(n_339), .B1(n_218), .B2(n_337), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_359), .B(n_339), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_364), .B(n_182), .C(n_200), .D(n_198), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_142), .B1(n_151), .B2(n_155), .C(n_237), .Y(n_398) );
OAI21xp33_ASAP7_75t_SL g399 ( .A1(n_365), .A2(n_150), .B(n_238), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_349), .A2(n_155), .B1(n_151), .B2(n_142), .C(n_303), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_396), .A2(n_155), .B(n_151), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
BUFx2_ASAP7_75t_SL g404 ( .A(n_376), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_373), .B(n_15), .C(n_16), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_371), .B(n_155), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_369), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_387), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_387), .B(n_150), .Y(n_412) );
AND2x4_ASAP7_75t_SL g413 ( .A(n_376), .B(n_337), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
INVxp33_ASAP7_75t_L g417 ( .A(n_368), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_383), .B(n_337), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_393), .B(n_15), .Y(n_419) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_373), .B(n_337), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_383), .B(n_337), .Y(n_421) );
AND2x2_ASAP7_75t_SL g422 ( .A(n_380), .B(n_272), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_384), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_390), .B(n_151), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_390), .B(n_16), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_375), .A2(n_139), .B1(n_272), .B2(n_273), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_393), .A2(n_18), .A3(n_194), .B1(n_185), .B2(n_183), .B3(n_260), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_372), .A2(n_398), .B(n_391), .Y(n_432) );
AOI33xp33_ASAP7_75t_L g433 ( .A1(n_383), .A2(n_194), .A3(n_18), .B1(n_260), .B2(n_215), .B3(n_253), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_377), .B(n_139), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
NOR2xp33_ASAP7_75t_R g436 ( .A(n_389), .B(n_273), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_229), .A3(n_279), .B(n_270), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_394), .B(n_273), .Y(n_439) );
AOI31xp33_ASAP7_75t_L g440 ( .A1(n_395), .A2(n_229), .A3(n_20), .B(n_21), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_394), .B(n_19), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_382), .Y(n_442) );
NAND3x1_ASAP7_75t_L g443 ( .A(n_400), .B(n_270), .C(n_293), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_382), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_399), .B(n_23), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_379), .B(n_273), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_378), .B(n_38), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_402), .Y(n_448) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_403), .A2(n_397), .A3(n_40), .B1(n_42), .B2(n_46), .B3(n_50), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_416), .B(n_39), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g451 ( .A(n_419), .B(n_272), .C(n_215), .D(n_270), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_415), .B(n_52), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_405), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_416), .B(n_54), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_427), .B(n_55), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_427), .B(n_56), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_415), .B(n_58), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_405), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_424), .B(n_61), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_248), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_417), .B(n_273), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_430), .B(n_251), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_425), .B(n_251), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_402), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_425), .B(n_248), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
INVxp33_ASAP7_75t_L g469 ( .A(n_436), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_414), .B(n_285), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_406), .B(n_287), .C(n_312), .D(n_297), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_408), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_413), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_414), .B(n_298), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_410), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_411), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_414), .B(n_287), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_404), .B(n_298), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_411), .B(n_298), .Y(n_480) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_404), .B(n_292), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_435), .B(n_297), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_428), .B(n_297), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_442), .B(n_252), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_433), .B(n_292), .C(n_191), .Y(n_488) );
NOR2x1p5_ASAP7_75t_L g489 ( .A(n_445), .B(n_312), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_401), .B(n_172), .C(n_191), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_420), .B(n_172), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_420), .B(n_293), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_413), .B(n_293), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_437), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_409), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_418), .B(n_253), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_418), .B(n_313), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_420), .B(n_172), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_482), .B(n_426), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_477), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_483), .B(n_426), .Y(n_501) );
NAND4xp75_ASAP7_75t_L g502 ( .A(n_491), .B(n_438), .C(n_422), .D(n_445), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_448), .B(n_442), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_453), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_491), .A2(n_440), .B(n_431), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_466), .B(n_444), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_472), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_448), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_487), .B(n_412), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_494), .B(n_444), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_495), .B(n_412), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_494), .B(n_437), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_474), .B(n_421), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_476), .B(n_421), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_456), .B(n_421), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_456), .B(n_465), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_473), .B(n_421), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_449), .A2(n_438), .B(n_447), .C(n_441), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g521 ( .A(n_462), .B(n_429), .C(n_447), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_486), .B(n_418), .Y(n_522) );
NAND3x1_ASAP7_75t_L g523 ( .A(n_481), .B(n_441), .C(n_446), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_451), .B(n_434), .C(n_439), .D(n_443), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_480), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_473), .B(n_413), .Y(n_526) );
AND4x1_ASAP7_75t_L g527 ( .A(n_488), .B(n_443), .C(n_422), .D(n_432), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g528 ( .A1(n_489), .A2(n_422), .A3(n_432), .B(n_197), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_470), .Y(n_529) );
NAND2x1p5_ASAP7_75t_SL g530 ( .A(n_479), .B(n_432), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_475), .B(n_172), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_464), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_469), .B(n_255), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_461), .B(n_191), .Y(n_534) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_469), .A2(n_191), .B(n_197), .Y(n_535) );
NAND4xp25_ASAP7_75t_L g536 ( .A(n_462), .B(n_210), .C(n_197), .D(n_212), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g537 ( .A1(n_471), .A2(n_197), .A3(n_210), .B(n_212), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_461), .B(n_210), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
OAI32xp33_ASAP7_75t_L g540 ( .A1(n_509), .A2(n_460), .A3(n_458), .B1(n_492), .B2(n_498), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_500), .B(n_463), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_532), .B(n_463), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_526), .B(n_450), .Y(n_543) );
NOR2xp67_ASAP7_75t_SL g544 ( .A(n_502), .B(n_536), .Y(n_544) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_526), .B(n_454), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_512), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_528), .A2(n_490), .B(n_454), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_539), .B(n_478), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_525), .B(n_478), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_505), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_512), .Y(n_552) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_518), .A2(n_450), .B(n_455), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_510), .Y(n_555) );
AOI21xp33_ASAP7_75t_L g556 ( .A1(n_520), .A2(n_457), .B(n_497), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_526), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_514), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_511), .B(n_484), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_503), .B(n_452), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_529), .B(n_485), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_527), .B(n_493), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_506), .A2(n_496), .B(n_217), .Y(n_563) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_523), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
XNOR2xp5_ASAP7_75t_L g566 ( .A(n_523), .B(n_217), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_508), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_508), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_521), .A2(n_217), .B(n_222), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_530), .A2(n_515), .B1(n_516), .B2(n_513), .C(n_501), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_522), .B(n_222), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g575 ( .A(n_524), .B(n_222), .Y(n_575) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_530), .B(n_534), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_533), .B(n_531), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_535), .A2(n_402), .B1(n_404), .B2(n_502), .Y(n_578) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_537), .B(n_538), .Y(n_579) );
XOR2xp5_ASAP7_75t_L g580 ( .A(n_519), .B(n_208), .Y(n_580) );
OAI211xp5_ASAP7_75t_SL g581 ( .A1(n_528), .A2(n_156), .B(n_80), .C(n_86), .Y(n_581) );
NOR3xp33_ASAP7_75t_SL g582 ( .A(n_528), .B(n_406), .C(n_502), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_509), .B(n_417), .Y(n_583) );
OAI31xp33_ASAP7_75t_L g584 ( .A1(n_564), .A2(n_578), .A3(n_562), .B(n_581), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_552), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_564), .A2(n_582), .B(n_556), .C(n_563), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_552), .Y(n_587) );
NAND3xp33_ASAP7_75t_SL g588 ( .A(n_578), .B(n_562), .C(n_571), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_555), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_583), .A2(n_570), .B(n_540), .C(n_568), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_545), .A2(n_557), .B1(n_543), .B2(n_558), .Y(n_591) );
AOI31xp33_ASAP7_75t_L g592 ( .A1(n_543), .A2(n_580), .A3(n_576), .B(n_547), .Y(n_592) );
OAI22x1_ASAP7_75t_L g593 ( .A1(n_558), .A2(n_566), .B1(n_560), .B2(n_551), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_567), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_542), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_592), .A2(n_572), .B1(n_559), .B2(n_548), .C(n_544), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_584), .A2(n_545), .B(n_579), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_586), .A2(n_559), .B(n_560), .C(n_546), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_588), .A2(n_570), .B(n_550), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_591), .A2(n_546), .B1(n_554), .B2(n_565), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_590), .A2(n_575), .B(n_553), .C(n_549), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_593), .A2(n_577), .B1(n_541), .B2(n_561), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_597), .A2(n_593), .B(n_594), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g604 ( .A1(n_598), .A2(n_585), .B(n_587), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_599), .B(n_595), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_602), .Y(n_606) );
AOI221xp5_ASAP7_75t_SL g607 ( .A1(n_603), .A2(n_596), .B1(n_600), .B2(n_601), .C(n_595), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_605), .A2(n_585), .B1(n_589), .B2(n_573), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_608), .B(n_606), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_607), .Y(n_610) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_610), .B(n_604), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_611), .B(n_609), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_612), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_613), .A2(n_574), .B(n_569), .Y(n_614) );
endmodule