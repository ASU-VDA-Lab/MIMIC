module fake_netlist_6_469_n_1939 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1939);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1939;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_8),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_45),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_95),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_19),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_59),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_114),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_105),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_136),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_40),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_3),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_75),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_132),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_124),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_115),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_184),
.Y(n_235)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_43),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_183),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_181),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_64),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_188),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_63),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_17),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_78),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_145),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_6),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_74),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_168),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_56),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_162),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_72),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_76),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_11),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_186),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_79),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_68),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_47),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_187),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_40),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_25),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_24),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_54),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_33),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_94),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_163),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_62),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_66),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_57),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_51),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_126),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_22),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_15),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_2),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_81),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_103),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_54),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_157),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_116),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_50),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_61),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_48),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_166),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_39),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_156),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_21),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_106),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_46),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_49),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_24),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_110),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_52),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_85),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_164),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_140),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_137),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_4),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_65),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_42),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_122),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_70),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_118),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_25),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_133),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_55),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_99),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_121),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_150),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_159),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_131),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_102),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_7),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_71),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_55),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_1),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_69),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_27),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_26),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_31),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_30),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_127),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_20),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_93),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_34),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_53),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_90),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_35),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_143),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_1),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_34),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_49),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_117),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_5),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_160),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_11),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_30),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_52),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_89),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_47),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_28),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_44),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_82),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_178),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_206),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_206),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_221),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_257),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_189),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_221),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_228),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_206),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_206),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_228),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_206),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_209),
.B(n_0),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_206),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_191),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_195),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_206),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_289),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_200),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_289),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_232),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_232),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_251),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_202),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_289),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_226),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_227),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_310),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_251),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_310),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_256),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_245),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_234),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_219),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_204),
.B(n_2),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_241),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_289),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_256),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_268),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_268),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_204),
.B(n_3),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_214),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_237),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_207),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_252),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_214),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_262),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_267),
.B(n_5),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_248),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_270),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_306),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_306),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_272),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_260),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_300),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_272),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_242),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_276),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_291),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_282),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_302),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_305),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_315),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_285),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_307),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_192),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_312),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_301),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_193),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_314),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_304),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_317),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_267),
.B(n_7),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_323),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_210),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_309),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_291),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_321),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_194),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_248),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_248),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_324),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_196),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_210),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_265),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_379),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_402),
.B(n_338),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_385),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_R g476 ( 
.A(n_394),
.B(n_295),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_451),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_386),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_378),
.B(n_231),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_454),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_415),
.B(n_376),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_421),
.B(n_197),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

NAND2x1_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_231),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_465),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_469),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_470),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_394),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_419),
.B(n_222),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_229),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

INVx6_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_395),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_384),
.B(n_244),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_420),
.B(n_222),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_395),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_375),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_398),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_422),
.B(n_357),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_425),
.B(n_241),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_390),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_384),
.B(n_299),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_398),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_413),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_430),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_413),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_460),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_408),
.B(n_203),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_470),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_424),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_424),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_231),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_438),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_470),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_442),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_404),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_426),
.B(n_243),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_410),
.B(n_208),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_463),
.Y(n_547)
);

AND3x1_ASAP7_75t_L g548 ( 
.A(n_392),
.B(n_344),
.C(n_339),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_463),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_503),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_503),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_504),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_486),
.B(n_412),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_483),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_519),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_510),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_486),
.B(n_407),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_509),
.B(n_406),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_516),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_485),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_522),
.B(n_229),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_490),
.B(n_249),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_490),
.B(n_442),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_514),
.B(n_445),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_407),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_441),
.B1(n_448),
.B2(n_414),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_528),
.B(n_380),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_528),
.B(n_445),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_548),
.B(n_249),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_370),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_480),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_516),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_453),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_480),
.B(n_449),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_533),
.A2(n_370),
.B1(n_354),
.B2(n_363),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_501),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_505),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_533),
.A2(n_372),
.B1(n_292),
.B2(n_434),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_516),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_501),
.B(n_449),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_546),
.B(n_456),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_546),
.B(n_231),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_533),
.B(n_456),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_473),
.B(n_190),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_505),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_550),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_550),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_502),
.B(n_461),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_483),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_487),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_516),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_521),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_502),
.B(n_461),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_502),
.B(n_464),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_383),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_505),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_533),
.B(n_214),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_541),
.B(n_466),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_508),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_533),
.A2(n_455),
.B1(n_446),
.B2(n_429),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_516),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_502),
.B(n_198),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_464),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_491),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_505),
.B(n_433),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_474),
.B(n_468),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_497),
.A2(n_381),
.B1(n_382),
.B2(n_468),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_416),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_508),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_491),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_507),
.A2(n_471),
.B1(n_443),
.B2(n_467),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_533),
.B(n_496),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_477),
.B(n_443),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_499),
.B(n_427),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_496),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_320),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_511),
.B(n_431),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_477),
.B(n_439),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_525),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_492),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_479),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_511),
.B(n_450),
.C(n_447),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_452),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_525),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_533),
.A2(n_459),
.B1(n_457),
.B2(n_318),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_481),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_473),
.B(n_199),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_481),
.B(n_488),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_265),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_513),
.A2(n_327),
.B1(n_374),
.B2(n_373),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_483),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_512),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_473),
.B(n_201),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_473),
.B(n_211),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_517),
.B(n_215),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_489),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_472),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_512),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_525),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_489),
.B(n_332),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_498),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_525),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_515),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_538),
.B(n_220),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_517),
.B(n_223),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_472),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_523),
.B(n_334),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_524),
.Y(n_672)
);

INVx8_ASAP7_75t_L g673 ( 
.A(n_483),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_525),
.B(n_212),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_475),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_518),
.B(n_238),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_492),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_482),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_498),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_512),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_540),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_500),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_540),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_483),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_483),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_526),
.B(n_347),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_495),
.Y(n_688)
);

BUFx4f_ASAP7_75t_L g689 ( 
.A(n_483),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_500),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_527),
.B(n_213),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_527),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_527),
.B(n_216),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_538),
.B(n_254),
.Y(n_697)
);

AND2x2_ASAP7_75t_SL g698 ( 
.A(n_518),
.B(n_273),
.Y(n_698)
);

AO22x2_ASAP7_75t_L g699 ( 
.A1(n_530),
.A2(n_293),
.B1(n_275),
.B2(n_279),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_540),
.A2(n_284),
.B1(n_325),
.B2(n_326),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_532),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_495),
.B(n_529),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_530),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_654),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_565),
.B(n_529),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_555),
.B(n_534),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_565),
.B(n_529),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_566),
.B(n_538),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_573),
.B(n_698),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_573),
.B(n_539),
.C(n_484),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_581),
.A2(n_205),
.B1(n_224),
.B2(n_230),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_569),
.A2(n_536),
.B(n_547),
.C(n_545),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_654),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_558),
.A2(n_341),
.B1(n_281),
.B2(n_294),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_348),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_601),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_L g717 ( 
.A(n_626),
.B(n_493),
.C(n_478),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_602),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_698),
.B(n_214),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_703),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_571),
.B(n_214),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_667),
.B(n_328),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_580),
.B(n_537),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_580),
.A2(n_389),
.B1(n_400),
.B2(n_401),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_675),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_572),
.B(n_214),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_596),
.B(n_599),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_660),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_575),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_596),
.B(n_537),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_599),
.A2(n_403),
.B1(n_409),
.B2(n_411),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_551),
.B(n_537),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_586),
.B(n_214),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_564),
.A2(n_333),
.B(n_340),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_595),
.B(n_322),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_579),
.B(n_350),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_670),
.B(n_610),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_553),
.B(n_346),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_554),
.B(n_542),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_557),
.B(n_542),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_562),
.B(n_542),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_661),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_563),
.B(n_549),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_575),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_570),
.B(n_549),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_570),
.B(n_549),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_651),
.B(n_494),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_621),
.B(n_217),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_665),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_671),
.B(n_356),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_585),
.B(n_218),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_359),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_648),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_656),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_600),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_625),
.B(n_225),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_662),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_625),
.B(n_361),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_688),
.B(n_535),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_581),
.B(n_233),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_582),
.B(n_535),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_603),
.B(n_362),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_634),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_690),
.B(n_322),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_672),
.Y(n_767)
);

BUFx2_ASAP7_75t_SL g768 ( 
.A(n_672),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_674),
.A2(n_547),
.B(n_545),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_637),
.B(n_568),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_659),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_582),
.B(n_536),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_603),
.B(n_367),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_582),
.B(n_543),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_582),
.A2(n_418),
.B1(n_436),
.B2(n_435),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_664),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_672),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_582),
.B(n_543),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_665),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_681),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_265),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_658),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_658),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_680),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_690),
.B(n_322),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_588),
.A2(n_239),
.B1(n_365),
.B2(n_352),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_588),
.A2(n_239),
.B1(n_365),
.B2(n_352),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_690),
.B(n_322),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_683),
.B(n_235),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_691),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_577),
.B(n_240),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_695),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_569),
.A2(n_290),
.B1(n_230),
.B2(n_224),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_702),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_694),
.B(n_246),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_552),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_583),
.B(n_250),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_587),
.B(n_255),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_687),
.B(n_368),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_598),
.B(n_685),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_590),
.B(n_258),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_608),
.B(n_371),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_593),
.B(n_259),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_650),
.B(n_261),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_650),
.B(n_263),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_592),
.A2(n_615),
.B1(n_700),
.B2(n_699),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_608),
.B(n_264),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_592),
.A2(n_366),
.B1(n_364),
.B2(n_360),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_693),
.B(n_269),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_696),
.B(n_277),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_679),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_616),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_658),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_627),
.B(n_278),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_682),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_609),
.B(n_280),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_685),
.B(n_322),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_627),
.B(n_283),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_633),
.B(n_313),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_552),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_685),
.B(n_322),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_600),
.Y(n_823)
);

INVx8_ASAP7_75t_L g824 ( 
.A(n_624),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_288),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_597),
.B(n_297),
.Y(n_826)
);

INVxp33_ASAP7_75t_L g827 ( 
.A(n_652),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_597),
.B(n_298),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_686),
.B(n_322),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_591),
.B(n_303),
.Y(n_830)
);

AND2x6_ASAP7_75t_SL g831 ( 
.A(n_676),
.B(n_205),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_609),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_591),
.B(n_308),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_682),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_556),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_701),
.B(n_313),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_311),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_686),
.B(n_632),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_615),
.A2(n_274),
.B1(n_290),
.B2(n_253),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_556),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_684),
.B(n_316),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_561),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_668),
.A2(n_358),
.B1(n_355),
.B2(n_353),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_692),
.B(n_319),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_335),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_663),
.A2(n_329),
.B(n_343),
.C(n_336),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_668),
.B(n_697),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_697),
.B(n_337),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_642),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_663),
.B(n_243),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_620),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_669),
.B(n_274),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_576),
.B(n_10),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_SL g854 ( 
.A(n_618),
.B(n_345),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_611),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_631),
.B(n_286),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_636),
.B(n_286),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_624),
.B(n_313),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_644),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_559),
.B(n_243),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_559),
.B(n_247),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_624),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_559),
.B(n_247),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_700),
.A2(n_345),
.B1(n_342),
.B2(n_253),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_611),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_567),
.B(n_247),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_686),
.B(n_330),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_561),
.Y(n_868)
);

BUFx5_ASAP7_75t_L g869 ( 
.A(n_620),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_574),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_673),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_669),
.A2(n_236),
.B1(n_287),
.B2(n_266),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_567),
.B(n_286),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_657),
.B(n_330),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_642),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_689),
.B(n_330),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_706),
.B(n_657),
.C(n_645),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_801),
.A2(n_689),
.B(n_673),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_801),
.A2(n_673),
.B(n_606),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_709),
.B(n_705),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_727),
.A2(n_647),
.B1(n_618),
.B2(n_678),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_838),
.A2(n_628),
.B(n_612),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_707),
.B(n_669),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_708),
.B(n_678),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_706),
.B(n_669),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_838),
.A2(n_673),
.B(n_641),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_816),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_760),
.A2(n_645),
.B(n_639),
.C(n_647),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_725),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_824),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_760),
.B(n_669),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_719),
.A2(n_622),
.B(n_612),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_770),
.B(n_676),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_SL g895 ( 
.A(n_871),
.B(n_560),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_723),
.A2(n_606),
.B(n_641),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_730),
.A2(n_606),
.B(n_641),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_871),
.A2(n_594),
.B(n_662),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_832),
.B(n_560),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_871),
.A2(n_594),
.B(n_662),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_727),
.A2(n_676),
.B1(n_677),
.B2(n_567),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_795),
.B(n_584),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_805),
.B(n_584),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_834),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_719),
.A2(n_622),
.B(n_628),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_808),
.B(n_560),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_806),
.B(n_584),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_871),
.A2(n_594),
.B(n_662),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_807),
.A2(n_677),
.B1(n_619),
.B2(n_646),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_720),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_763),
.A2(n_774),
.B(n_772),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_766),
.A2(n_614),
.B(n_630),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_778),
.A2(n_666),
.B(n_640),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_759),
.A2(n_666),
.B(n_640),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_766),
.A2(n_613),
.B(n_623),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_761),
.A2(n_666),
.B(n_604),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_867),
.A2(n_666),
.B(n_604),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_867),
.A2(n_560),
.B(n_604),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_810),
.A2(n_640),
.B(n_604),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_797),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_807),
.A2(n_677),
.B1(n_619),
.B2(n_646),
.Y(n_921)
);

AO22x1_ASAP7_75t_L g922 ( 
.A1(n_827),
.A2(n_655),
.B1(n_649),
.B2(n_620),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_821),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_808),
.B(n_640),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_820),
.B(n_646),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_745),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_755),
.B(n_619),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_817),
.B(n_653),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_728),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_738),
.B(n_266),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_811),
.A2(n_653),
.B(n_578),
.Y(n_931)
);

AO21x1_ASAP7_75t_L g932 ( 
.A1(n_734),
.A2(n_605),
.B(n_638),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_756),
.B(n_771),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_L g934 ( 
.A(n_767),
.B(n_639),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_734),
.A2(n_574),
.B(n_578),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_769),
.A2(n_748),
.B(n_747),
.Y(n_936)
);

AO21x1_ASAP7_75t_L g937 ( 
.A1(n_736),
.A2(n_635),
.B(n_629),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_837),
.A2(n_653),
.B(n_617),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_875),
.B(n_653),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_754),
.B(n_287),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_764),
.A2(n_629),
.B(n_635),
.C(n_617),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_736),
.A2(n_699),
.B(n_620),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_812),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_813),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_817),
.B(n_342),
.Y(n_946)
);

NOR2x1_ASAP7_75t_L g947 ( 
.A(n_768),
.B(n_699),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_784),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_841),
.A2(n_620),
.B(n_655),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_781),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_836),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_844),
.A2(n_845),
.B(n_833),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_791),
.B(n_655),
.Y(n_953)
);

NOR2x1_ASAP7_75t_L g954 ( 
.A(n_749),
.B(n_655),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_830),
.A2(n_655),
.B(n_649),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_716),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_718),
.B(n_649),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_818),
.A2(n_829),
.B(n_822),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_754),
.B(n_649),
.C(n_12),
.Y(n_959)
);

OA22x2_ASAP7_75t_L g960 ( 
.A1(n_864),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_818),
.A2(n_649),
.B(n_88),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_822),
.A2(n_87),
.B(n_177),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_850),
.B(n_13),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_829),
.A2(n_84),
.B(n_176),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_875),
.B(n_80),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_792),
.A2(n_92),
.B(n_175),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_777),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_793),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_835),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_815),
.B(n_14),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_798),
.A2(n_77),
.B(n_167),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_782),
.B(n_67),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_799),
.A2(n_96),
.B(n_158),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_783),
.A2(n_60),
.B1(n_154),
.B2(n_147),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_802),
.A2(n_182),
.B(n_138),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_840),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_762),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_819),
.B(n_16),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_804),
.A2(n_135),
.B(n_134),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_129),
.B(n_125),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_785),
.A2(n_120),
.B(n_112),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_788),
.A2(n_100),
.B(n_98),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_788),
.A2(n_97),
.B(n_27),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_847),
.A2(n_714),
.B(n_794),
.C(n_876),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_825),
.B(n_23),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_737),
.B(n_23),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_765),
.B(n_29),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_737),
.B(n_32),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_721),
.A2(n_726),
.B(n_733),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_729),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_721),
.A2(n_32),
.B(n_38),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_764),
.A2(n_56),
.B(n_41),
.C(n_44),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_726),
.A2(n_38),
.B(n_41),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_852),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_824),
.B(n_722),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_814),
.A2(n_744),
.B(n_741),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_859),
.A2(n_870),
.B(n_842),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_773),
.A2(n_803),
.B(n_876),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_773),
.B(n_803),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_872),
.B(n_849),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_868),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_874),
.B(n_854),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_746),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_740),
.A2(n_742),
.B(n_729),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_874),
.A2(n_715),
.B(n_858),
.C(n_712),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_704),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_786),
.B(n_787),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_846),
.A2(n_743),
.B(n_780),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_715),
.B(n_758),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_713),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_729),
.A2(n_855),
.B(n_865),
.Y(n_1011)
);

CKINVDCx8_ASAP7_75t_R g1012 ( 
.A(n_831),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_724),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_752),
.B(n_800),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_731),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_786),
.A2(n_787),
.B(n_839),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_862),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_739),
.B(n_823),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_839),
.A2(n_823),
.B1(n_757),
.B2(n_865),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_757),
.B(n_789),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_794),
.A2(n_809),
.B(n_858),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_729),
.A2(n_855),
.B(n_751),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_779),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_790),
.A2(n_828),
.B(n_826),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_860),
.A2(n_873),
.B(n_866),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_861),
.Y(n_1026)
);

INVx3_ASAP7_75t_SL g1027 ( 
.A(n_722),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_863),
.A2(n_735),
.B(n_857),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_775),
.B(n_732),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_824),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_853),
.Y(n_1031)
);

NAND2x1_ASAP7_75t_L g1032 ( 
.A(n_851),
.B(n_869),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_753),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_796),
.B(n_722),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_848),
.A2(n_750),
.B(n_856),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_843),
.A2(n_710),
.B(n_717),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_851),
.A2(n_869),
.B(n_711),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_851),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_711),
.B(n_851),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_851),
.B(n_869),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_851),
.A2(n_801),
.B(n_838),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_869),
.A2(n_709),
.B1(n_727),
.B2(n_807),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_869),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_869),
.B(n_709),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_709),
.B(n_705),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_816),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_770),
.B(n_566),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_709),
.B(n_708),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_709),
.B(n_708),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_709),
.A2(n_569),
.B(n_727),
.C(n_760),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_816),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_816),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_709),
.B(n_705),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1061)
);

NOR2x1p5_ASAP7_75t_L g1062 ( 
.A(n_767),
.B(n_478),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_760),
.A2(n_709),
.B(n_565),
.C(n_573),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_801),
.A2(n_838),
.B(n_730),
.Y(n_1064)
);

AO22x1_ASAP7_75t_L g1065 ( 
.A1(n_760),
.A2(n_827),
.B1(n_709),
.B2(n_706),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_709),
.A2(n_727),
.B1(n_807),
.B2(n_832),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_746),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_709),
.B(n_708),
.Y(n_1068)
);

OAI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_709),
.A2(n_827),
.B1(n_832),
.B2(n_727),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_709),
.A2(n_569),
.B(n_727),
.C(n_760),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_911),
.A2(n_958),
.B(n_1025),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_999),
.B(n_1063),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_1016),
.B(n_1007),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_929),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_944),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_881),
.B(n_1045),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1047),
.A2(n_1052),
.B(n_1049),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_910),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_984),
.A2(n_1021),
.B(n_941),
.C(n_1070),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_926),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_938),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_935),
.A2(n_936),
.B(n_883),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_SL g1084 ( 
.A(n_1030),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_1030),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1060),
.B(n_1065),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1047),
.A2(n_1052),
.B(n_1049),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_890),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1042),
.A2(n_1057),
.B(n_1053),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1057),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1030),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1054),
.A2(n_1039),
.B(n_988),
.C(n_986),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1004),
.A2(n_989),
.B(n_879),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1048),
.B(n_930),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1058),
.A2(n_1061),
.B(n_1059),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1003),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_967),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1059),
.A2(n_1064),
.B(n_1061),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1068),
.B(n_1069),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_948),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1013),
.A2(n_1014),
.B1(n_1036),
.B2(n_1009),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_995),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1064),
.A2(n_892),
.B(n_886),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1003),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_889),
.A2(n_1066),
.B1(n_1002),
.B2(n_946),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_998),
.A2(n_877),
.B1(n_1000),
.B2(n_963),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_989),
.A2(n_879),
.B(n_893),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1017),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_891),
.B(n_1003),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_945),
.B(n_1031),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1005),
.A2(n_1035),
.B(n_1037),
.C(n_970),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_995),
.B(n_1067),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_950),
.B(n_951),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_894),
.B(n_934),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_978),
.A2(n_985),
.B(n_1033),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_906),
.A2(n_928),
.B(n_924),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1026),
.B(n_933),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1020),
.B(n_885),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_956),
.B(n_1018),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_905),
.A2(n_1032),
.B(n_896),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_884),
.A2(n_1044),
.B(n_1028),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_968),
.B(n_880),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1067),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_953),
.A2(n_957),
.B(n_925),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_880),
.B(n_1035),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_SL g1127 ( 
.A1(n_972),
.A2(n_902),
.B(n_907),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_932),
.A2(n_937),
.A3(n_942),
.B(n_901),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_995),
.B(n_1067),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_909),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_972),
.B(n_997),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_994),
.B(n_977),
.C(n_992),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_896),
.A2(n_897),
.B(n_887),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1041),
.A2(n_887),
.B(n_952),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_959),
.B(n_1029),
.C(n_987),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_891),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1037),
.A2(n_882),
.B(n_1041),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_903),
.A2(n_878),
.B(n_897),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1028),
.A2(n_943),
.B(n_996),
.C(n_1024),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_943),
.A2(n_962),
.B(n_947),
.C(n_1034),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1046),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1142)
);

AOI221xp5_ASAP7_75t_L g1143 ( 
.A1(n_991),
.A2(n_993),
.B1(n_974),
.B2(n_1056),
.C(n_1055),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_990),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_898),
.A2(n_900),
.B(n_908),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1012),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_878),
.A2(n_1040),
.B(n_949),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1062),
.B(n_960),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_954),
.B(n_990),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_888),
.B(n_923),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_1008),
.A2(n_955),
.B(n_921),
.Y(n_1151)
);

NAND2x1_ASAP7_75t_L g1152 ( 
.A(n_895),
.B(n_1043),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_960),
.A2(n_927),
.B1(n_1038),
.B2(n_1015),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_920),
.B(n_969),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_961),
.A2(n_983),
.A3(n_917),
.B(n_973),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_976),
.B(n_1001),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1006),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1023),
.B(n_1010),
.Y(n_1158)
);

BUFx4f_ASAP7_75t_SL g1159 ( 
.A(n_965),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1011),
.A2(n_1022),
.B(n_913),
.Y(n_1160)
);

AOI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_899),
.A2(n_940),
.B(n_931),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_922),
.B(n_940),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_916),
.A2(n_914),
.B(n_939),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_918),
.A2(n_919),
.B(n_964),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_980),
.B(n_981),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_982),
.A2(n_966),
.B(n_971),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_975),
.A2(n_979),
.B(n_999),
.C(n_1063),
.Y(n_1167)
);

AND3x2_ASAP7_75t_L g1168 ( 
.A(n_1007),
.B(n_999),
.C(n_941),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_929),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_911),
.A2(n_871),
.B(n_801),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_999),
.A2(n_1063),
.B1(n_709),
.B2(n_1016),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_999),
.A2(n_1063),
.B(n_984),
.C(n_709),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_929),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_999),
.B(n_1063),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_990),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_944),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_SL g1178 ( 
.A(n_1016),
.B(n_999),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_998),
.A2(n_932),
.A3(n_1042),
.B(n_937),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_999),
.B(n_832),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_999),
.A2(n_1063),
.B(n_998),
.C(n_1065),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_999),
.B(n_1063),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_944),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1048),
.B(n_708),
.Y(n_1184)
);

OAI21xp33_ASAP7_75t_SL g1185 ( 
.A1(n_999),
.A2(n_807),
.B(n_1002),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_998),
.A2(n_932),
.A3(n_1042),
.B(n_937),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_999),
.A2(n_1042),
.B(n_1063),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_999),
.B(n_1063),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_999),
.B(n_1063),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_999),
.A2(n_1063),
.B(n_984),
.C(n_709),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_999),
.A2(n_941),
.B(n_709),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_999),
.A2(n_941),
.B(n_709),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_SL g1195 ( 
.A1(n_999),
.A2(n_807),
.B(n_1002),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_999),
.A2(n_1063),
.B(n_984),
.C(n_709),
.Y(n_1196)
);

OA22x2_ASAP7_75t_L g1197 ( 
.A1(n_1016),
.A2(n_1007),
.B1(n_864),
.B2(n_946),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_910),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_999),
.B(n_1063),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1030),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1030),
.B(n_891),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_911),
.A2(n_871),
.B(n_801),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_999),
.A2(n_709),
.B1(n_941),
.B2(n_986),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_911),
.A2(n_871),
.B(n_801),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_999),
.B(n_1063),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_990),
.Y(n_1207)
);

AND2x2_ASAP7_75t_SL g1208 ( 
.A(n_1007),
.B(n_999),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_998),
.A2(n_932),
.A3(n_1042),
.B(n_937),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_999),
.A2(n_1039),
.B1(n_1063),
.B2(n_709),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_999),
.A2(n_1063),
.B(n_984),
.C(n_709),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1048),
.B(n_708),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_911),
.A2(n_871),
.B(n_801),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_906),
.A2(n_928),
.B(n_924),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_999),
.A2(n_1063),
.B1(n_709),
.B2(n_1039),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_999),
.B(n_1063),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_911),
.A2(n_871),
.B(n_801),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_SL g1219 ( 
.A1(n_999),
.A2(n_1042),
.B(n_1044),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_L g1220 ( 
.A(n_1062),
.B(n_768),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_999),
.A2(n_1042),
.B(n_1063),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_935),
.A2(n_915),
.B(n_912),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_999),
.A2(n_1042),
.B(n_1044),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1030),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_998),
.A2(n_932),
.A3(n_1042),
.B(n_937),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_904),
.Y(n_1226)
);

AOI21xp33_ASAP7_75t_L g1227 ( 
.A1(n_999),
.A2(n_941),
.B(n_709),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_999),
.A2(n_1042),
.B(n_1063),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_999),
.B(n_1063),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_999),
.B(n_1044),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1076),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1193),
.B(n_1194),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1078),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1081),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1227),
.A2(n_1079),
.B(n_1185),
.C(n_1195),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1203),
.A2(n_1116),
.B(n_1196),
.C(n_1211),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1082),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1103),
.B(n_1136),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1075),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1102),
.B(n_1184),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1094),
.B(n_1212),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1101),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1198),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1103),
.B(n_1136),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

AO21x2_ASAP7_75t_L g1246 ( 
.A1(n_1090),
.A2(n_1089),
.B(n_1087),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1144),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1074),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1187),
.A2(n_1228),
.B(n_1221),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1197),
.A2(n_1208),
.B1(n_1178),
.B2(n_1106),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1091),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1103),
.B(n_1113),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1089),
.A2(n_1090),
.B(n_1112),
.Y(n_1253)
);

CKINVDCx8_ASAP7_75t_R g1254 ( 
.A(n_1088),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1115),
.B(n_1111),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1109),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1177),
.B(n_1183),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1169),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1142),
.B(n_1148),
.Y(n_1259)
);

O2A1O1Ixp5_ASAP7_75t_SL g1260 ( 
.A1(n_1106),
.A2(n_1171),
.B(n_1216),
.C(n_1187),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1118),
.B(n_1086),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1113),
.B(n_1129),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1173),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1178),
.A2(n_1221),
.B1(n_1228),
.B2(n_1135),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1091),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1144),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1124),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1113),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1129),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1114),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1129),
.B(n_1085),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1201),
.B(n_1110),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1172),
.A2(n_1192),
.B(n_1185),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1210),
.A2(n_1182),
.B1(n_1199),
.B2(n_1072),
.Y(n_1274)
);

O2A1O1Ixp5_ASAP7_75t_L g1275 ( 
.A1(n_1167),
.A2(n_1181),
.B(n_1166),
.C(n_1092),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1098),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1120),
.B(n_1180),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1175),
.B(n_1189),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1071),
.A2(n_1202),
.B(n_1213),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1146),
.Y(n_1280)
);

O2A1O1Ixp5_ASAP7_75t_L g1281 ( 
.A1(n_1171),
.A2(n_1217),
.B(n_1229),
.C(n_1206),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1134),
.A2(n_1104),
.B(n_1139),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1191),
.B(n_1210),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1144),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1170),
.A2(n_1205),
.B(n_1218),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1195),
.A2(n_1100),
.B(n_1140),
.C(n_1131),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1219),
.A2(n_1223),
.B(n_1165),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1130),
.B(n_1073),
.Y(n_1288)
);

O2A1O1Ixp5_ASAP7_75t_L g1289 ( 
.A1(n_1163),
.A2(n_1077),
.B(n_1099),
.C(n_1095),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1138),
.A2(n_1137),
.B(n_1160),
.Y(n_1290)
);

O2A1O1Ixp5_ASAP7_75t_L g1291 ( 
.A1(n_1147),
.A2(n_1122),
.B(n_1132),
.C(n_1161),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1073),
.B(n_1230),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1180),
.B(n_1226),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1159),
.A2(n_1132),
.B1(n_1135),
.B2(n_1084),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1141),
.B(n_1150),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1151),
.A2(n_1126),
.B(n_1133),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1230),
.B(n_1096),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1151),
.A2(n_1093),
.B(n_1108),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1084),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1085),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1230),
.B(n_1119),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1176),
.B(n_1207),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1168),
.B(n_1097),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1097),
.B(n_1105),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1230),
.A2(n_1107),
.B1(n_1153),
.B2(n_1143),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1091),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1154),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1123),
.A2(n_1153),
.B1(n_1156),
.B2(n_1158),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1149),
.B(n_1179),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1200),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1097),
.Y(n_1312)
);

BUFx2_ASAP7_75t_R g1313 ( 
.A(n_1162),
.Y(n_1313)
);

BUFx8_ASAP7_75t_L g1314 ( 
.A(n_1200),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1149),
.B(n_1179),
.Y(n_1315)
);

INVx5_ASAP7_75t_L g1316 ( 
.A(n_1200),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1224),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1105),
.B(n_1224),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1220),
.A2(n_1207),
.B(n_1152),
.C(n_1127),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1121),
.A2(n_1145),
.B(n_1164),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1224),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1117),
.A2(n_1215),
.B1(n_1186),
.B2(n_1225),
.Y(n_1322)
);

O2A1O1Ixp5_ASAP7_75t_SL g1323 ( 
.A1(n_1125),
.A2(n_1225),
.B(n_1209),
.C(n_1186),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1080),
.B(n_1190),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1209),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1209),
.B(n_1225),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1083),
.A2(n_1188),
.B(n_1222),
.Y(n_1327)
);

CKINVDCx8_ASAP7_75t_R g1328 ( 
.A(n_1128),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1174),
.B(n_1204),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1155),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1128),
.B(n_1214),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1155),
.B(n_1076),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1155),
.B(n_1076),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1074),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1094),
.B(n_1048),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1075),
.B(n_738),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1103),
.B(n_1136),
.Y(n_1337)
);

INVx3_ASAP7_75t_R g1338 ( 
.A(n_1088),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1074),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1136),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1076),
.B(n_999),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1094),
.B(n_1048),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1103),
.B(n_1136),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1088),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1094),
.B(n_1048),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1075),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1193),
.A2(n_1063),
.B(n_999),
.C(n_1227),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1074),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1071),
.A2(n_1202),
.B(n_1170),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1193),
.A2(n_1063),
.B(n_999),
.C(n_1227),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1076),
.A2(n_999),
.B1(n_1063),
.B2(n_1016),
.Y(n_1351)
);

INVx5_ASAP7_75t_L g1352 ( 
.A(n_1144),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1193),
.A2(n_999),
.B(n_1063),
.C(n_1227),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1074),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1170),
.A2(n_1205),
.B(n_1202),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1075),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1075),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1203),
.A2(n_999),
.B1(n_941),
.B2(n_1016),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1078),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1088),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1076),
.A2(n_999),
.B1(n_1063),
.B2(n_1016),
.Y(n_1361)
);

OA22x2_ASAP7_75t_L g1362 ( 
.A1(n_1094),
.A2(n_1016),
.B1(n_1007),
.B2(n_946),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1103),
.B(n_1136),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1094),
.B(n_1048),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1075),
.B(n_738),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1076),
.A2(n_999),
.B1(n_1063),
.B2(n_1016),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1113),
.B(n_768),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1076),
.B(n_999),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1071),
.A2(n_1202),
.B(n_1170),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1078),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1136),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1178),
.A2(n_999),
.B1(n_709),
.B2(n_941),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1076),
.B(n_999),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1074),
.Y(n_1374)
);

INVx2_ASAP7_75t_R g1375 ( 
.A(n_1103),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1203),
.A2(n_999),
.B1(n_941),
.B2(n_1016),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1111),
.Y(n_1377)
);

OR2x6_ASAP7_75t_SL g1378 ( 
.A(n_1135),
.B(n_478),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1102),
.B(n_999),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1379),
.A2(n_1358),
.B1(n_1376),
.B2(n_1249),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1338),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1257),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1358),
.A2(n_1376),
.B1(n_1249),
.B2(n_1372),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1356),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1275),
.A2(n_1282),
.B(n_1289),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1327),
.A2(n_1287),
.B(n_1296),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1241),
.B(n_1335),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1237),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1280),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1242),
.Y(n_1390)
);

INVx3_ASAP7_75t_SL g1391 ( 
.A(n_1276),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1243),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1247),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1240),
.B(n_1341),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1341),
.B(n_1368),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1353),
.A2(n_1350),
.B(n_1347),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1239),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1346),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1357),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1247),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1254),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1368),
.A2(n_1373),
.B1(n_1255),
.B2(n_1273),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1370),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1247),
.B(n_1352),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1234),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1264),
.A2(n_1232),
.B1(n_1250),
.B2(n_1366),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1290),
.A2(n_1279),
.B(n_1369),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1373),
.A2(n_1231),
.B1(n_1377),
.B2(n_1294),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1314),
.Y(n_1409)
);

CKINVDCx6p67_ASAP7_75t_R g1410 ( 
.A(n_1352),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1261),
.B(n_1342),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1352),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1316),
.Y(n_1413)
);

AO21x1_ASAP7_75t_L g1414 ( 
.A1(n_1236),
.A2(n_1351),
.B(n_1361),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_R g1415 ( 
.A1(n_1270),
.A2(n_1336),
.B1(n_1365),
.B2(n_1256),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_L g1416 ( 
.A1(n_1232),
.A2(n_1235),
.B(n_1306),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1351),
.A2(n_1361),
.B1(n_1366),
.B2(n_1362),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1378),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1274),
.A2(n_1286),
.B(n_1302),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1344),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1303),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1274),
.A2(n_1302),
.B(n_1306),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1270),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1359),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1248),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1267),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1316),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1345),
.B(n_1364),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1314),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1320),
.A2(n_1355),
.B(n_1298),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1295),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1273),
.A2(n_1259),
.B1(n_1362),
.B2(n_1277),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1324),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1301),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1308),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1293),
.B(n_1304),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1262),
.B(n_1268),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1246),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1283),
.A2(n_1252),
.B1(n_1253),
.B2(n_1360),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1246),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1283),
.A2(n_1278),
.B1(n_1313),
.B2(n_1288),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1310),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1288),
.Y(n_1444)
);

NOR2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1334),
.B(n_1348),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1278),
.A2(n_1253),
.B1(n_1309),
.B2(n_1297),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1367),
.A2(n_1292),
.B1(n_1297),
.B2(n_1271),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1324),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1329),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1307),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1263),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1245),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1310),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1266),
.Y(n_1454)
);

INVxp33_ASAP7_75t_L g1455 ( 
.A(n_1312),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1271),
.B(n_1238),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1238),
.B(n_1244),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1315),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1339),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1329),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1324),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1354),
.Y(n_1463)
);

CKINVDCx8_ASAP7_75t_R g1464 ( 
.A(n_1300),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1374),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1272),
.B(n_1367),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1305),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1245),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1292),
.A2(n_1244),
.B1(n_1337),
.B2(n_1343),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1309),
.A2(n_1333),
.B1(n_1332),
.B2(n_1330),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1245),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1285),
.A2(n_1296),
.B(n_1282),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1332),
.B(n_1333),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1315),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1326),
.A2(n_1325),
.B1(n_1375),
.B2(n_1272),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1272),
.B(n_1313),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1340),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1337),
.A2(n_1363),
.B1(n_1343),
.B2(n_1371),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1305),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1266),
.B(n_1284),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1363),
.B(n_1284),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1319),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1322),
.A2(n_1331),
.B1(n_1299),
.B2(n_1318),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1251),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1291),
.Y(n_1485)
);

BUFx2_ASAP7_75t_R g1486 ( 
.A(n_1328),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1322),
.A2(n_1317),
.B1(n_1311),
.B2(n_1251),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1281),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1265),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1349),
.A2(n_1323),
.B(n_1321),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1314),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1280),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1254),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1379),
.A2(n_999),
.B1(n_941),
.B2(n_385),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1241),
.B(n_1335),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1247),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1257),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1233),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1233),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1252),
.B(n_1262),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1254),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1231),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1303),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1356),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1379),
.A2(n_999),
.B1(n_1368),
.B2(n_1341),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1443),
.B(n_1453),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1502),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1433),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1386),
.A2(n_1430),
.B(n_1407),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1458),
.B(n_1474),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1396),
.B(n_1473),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1423),
.Y(n_1513)
);

BUFx2_ASAP7_75t_SL g1514 ( 
.A(n_1464),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1444),
.B(n_1380),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1380),
.B(n_1417),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1433),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1430),
.A2(n_1488),
.B(n_1470),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1439),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1414),
.A2(n_1472),
.B(n_1490),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1485),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1417),
.B(n_1416),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1462),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1433),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1422),
.B(n_1406),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1406),
.B(n_1470),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1485),
.A2(n_1446),
.B(n_1419),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1441),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1384),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1446),
.B(n_1394),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1448),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1385),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1385),
.A2(n_1449),
.B(n_1461),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

AO21x1_ASAP7_75t_SL g1535 ( 
.A1(n_1383),
.A2(n_1475),
.B(n_1460),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1427),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1472),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1408),
.B(n_1505),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1482),
.A2(n_1394),
.B(n_1405),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1432),
.B(n_1402),
.Y(n_1540)
);

INVx8_ASAP7_75t_L g1541 ( 
.A(n_1427),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1424),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1383),
.A2(n_1494),
.B(n_1395),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1431),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1411),
.B(n_1483),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1475),
.A2(n_1483),
.B(n_1421),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1395),
.B(n_1390),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1435),
.Y(n_1549)
);

BUFx2_ASAP7_75t_R g1550 ( 
.A(n_1409),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1397),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1388),
.Y(n_1552)
);

OR2x6_ASAP7_75t_L g1553 ( 
.A(n_1427),
.B(n_1421),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1392),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1442),
.A2(n_1498),
.B(n_1403),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1382),
.B(n_1497),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1503),
.B(n_1500),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1387),
.B(n_1495),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1456),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1499),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1398),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1447),
.B(n_1440),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1426),
.Y(n_1563)
);

NAND2x1p5_ASAP7_75t_L g1564 ( 
.A(n_1413),
.B(n_1496),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1493),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1434),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1487),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1428),
.B(n_1500),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1393),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1393),
.Y(n_1570)
);

BUFx12f_ASAP7_75t_L g1571 ( 
.A(n_1493),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1479),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1500),
.B(n_1436),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1454),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1399),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1489),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1480),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1404),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1481),
.B(n_1457),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1418),
.B(n_1469),
.C(n_1463),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1455),
.A2(n_1478),
.B(n_1457),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1415),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1457),
.B(n_1467),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1486),
.B(n_1476),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1518),
.B(n_1455),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1544),
.A2(n_1418),
.B1(n_1451),
.B2(n_1381),
.Y(n_1587)
);

AND2x4_ASAP7_75t_SL g1588 ( 
.A(n_1553),
.B(n_1410),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1539),
.B(n_1465),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1518),
.B(n_1484),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1521),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1544),
.A2(n_1381),
.B1(n_1391),
.B2(n_1420),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1539),
.B(n_1391),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1539),
.B(n_1459),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1389),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1512),
.B(n_1400),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1528),
.B(n_1520),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1532),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1512),
.B(n_1412),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_SL g1601 ( 
.A(n_1535),
.B(n_1412),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1507),
.B(n_1515),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1520),
.B(n_1452),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1521),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1533),
.B(n_1539),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1561),
.Y(n_1607)
);

OA21x2_ASAP7_75t_L g1608 ( 
.A1(n_1510),
.A2(n_1468),
.B(n_1425),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1507),
.B(n_1412),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1515),
.B(n_1412),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1538),
.A2(n_1401),
.B(n_1468),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1527),
.B(n_1471),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1527),
.B(n_1523),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1526),
.A2(n_1401),
.B1(n_1491),
.B2(n_1409),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1527),
.B(n_1471),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1527),
.B(n_1429),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1534),
.B(n_1429),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1561),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1511),
.B(n_1530),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1549),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1524),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1513),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1553),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1545),
.B(n_1548),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1593),
.A2(n_1581),
.B(n_1538),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1606),
.A2(n_1510),
.B(n_1537),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1617),
.B(n_1509),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1594),
.B(n_1525),
.C(n_1583),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1601),
.A2(n_1525),
.B(n_1581),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1624),
.B(n_1627),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1627),
.B(n_1583),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1611),
.B(n_1562),
.C(n_1582),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1621),
.B(n_1513),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1615),
.B(n_1557),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1587),
.A2(n_1540),
.B(n_1526),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1621),
.B(n_1545),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1617),
.B(n_1618),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1618),
.B(n_1509),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_SL g1642 ( 
.A(n_1611),
.B(n_1540),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1548),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1618),
.B(n_1625),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_L g1645 ( 
.A(n_1594),
.B(n_1546),
.C(n_1556),
.D(n_1529),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1615),
.A2(n_1522),
.B(n_1562),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1596),
.A2(n_1522),
.B(n_1516),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1625),
.B(n_1508),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1620),
.B(n_1529),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1606),
.A2(n_1510),
.B(n_1589),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1597),
.A2(n_1550),
.B1(n_1546),
.B2(n_1516),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1602),
.B(n_1543),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1625),
.B(n_1508),
.Y(n_1653)
);

NAND4xp25_ASAP7_75t_L g1654 ( 
.A(n_1590),
.B(n_1543),
.C(n_1567),
.D(n_1558),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1577),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1508),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1599),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1586),
.B(n_1517),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1590),
.A2(n_1567),
.B(n_1550),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1586),
.B(n_1517),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1600),
.B(n_1577),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1600),
.A2(n_1514),
.B1(n_1610),
.B2(n_1582),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1626),
.A2(n_1535),
.B1(n_1555),
.B2(n_1557),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1610),
.B(n_1558),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1609),
.B(n_1551),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1609),
.B(n_1563),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_SL g1669 ( 
.A1(n_1612),
.A2(n_1547),
.B(n_1574),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1595),
.A2(n_1575),
.B1(n_1549),
.B2(n_1552),
.C(n_1576),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1595),
.B(n_1542),
.C(n_1560),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1588),
.A2(n_1585),
.B(n_1573),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1612),
.B(n_1542),
.C(n_1560),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1622),
.A2(n_1552),
.B1(n_1576),
.B2(n_1554),
.C(n_1566),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1622),
.A2(n_1554),
.B1(n_1566),
.B2(n_1578),
.C(n_1555),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1612),
.B(n_1574),
.C(n_1572),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1614),
.B(n_1555),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1616),
.A2(n_1585),
.B1(n_1568),
.B2(n_1573),
.C(n_1578),
.Y(n_1679)
);

OAI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1616),
.A2(n_1568),
.B(n_1547),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1616),
.B(n_1572),
.C(n_1579),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1619),
.B(n_1555),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1603),
.B(n_1531),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1659),
.Y(n_1684)
);

INVx5_ASAP7_75t_L g1685 ( 
.A(n_1659),
.Y(n_1685)
);

INVx5_ASAP7_75t_L g1686 ( 
.A(n_1660),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1678),
.B(n_1613),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1682),
.B(n_1613),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1642),
.A2(n_1514),
.B1(n_1580),
.B2(n_1584),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1662),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1639),
.B(n_1605),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1605),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1650),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1628),
.A2(n_1626),
.B1(n_1553),
.B2(n_1559),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1592),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1642),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1634),
.B(n_1598),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1640),
.B(n_1644),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1650),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1631),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1650),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1630),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1683),
.B(n_1680),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1571),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1629),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1680),
.B(n_1591),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1598),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1636),
.B(n_1598),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1629),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1681),
.B(n_1626),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1657),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1686),
.B(n_1674),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1658),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1668),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1706),
.B(n_1648),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1703),
.B(n_1666),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1685),
.B(n_1608),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1686),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1709),
.A2(n_1647),
.B1(n_1638),
.B2(n_1635),
.C(n_1646),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1715),
.B(n_1632),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1706),
.B(n_1648),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

AND2x4_ASAP7_75t_SL g1731 ( 
.A(n_1691),
.B(n_1641),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1684),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1708),
.B(n_1643),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1710),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1707),
.B(n_1571),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1710),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1649),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1698),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1715),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1687),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1714),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1686),
.B(n_1626),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1716),
.B(n_1654),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1698),
.B(n_1653),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1693),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1713),
.B(n_1641),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1689),
.B(n_1671),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1632),
.Y(n_1752)
);

NAND4xp25_ASAP7_75t_L g1753 ( 
.A(n_1712),
.B(n_1665),
.C(n_1661),
.D(n_1679),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1656),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1695),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1726),
.B(n_1711),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1751),
.B(n_1712),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1742),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1735),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1741),
.B(n_1711),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1741),
.B(n_1701),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1745),
.Y(n_1762)
);

AND2x2_ASAP7_75t_SL g1763 ( 
.A(n_1717),
.B(n_1731),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1728),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1742),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1722),
.A2(n_1699),
.B1(n_1691),
.B2(n_1728),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1735),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1755),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1725),
.B(n_1700),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1752),
.B(n_1701),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1752),
.B(n_1705),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1746),
.B(n_1700),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1724),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1747),
.B(n_1690),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1739),
.B(n_1690),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1753),
.B(n_1661),
.C(n_1651),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1740),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1751),
.B(n_1713),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1749),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1718),
.B(n_1695),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1738),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_SL g1784 ( 
.A1(n_1731),
.A2(n_1601),
.B1(n_1686),
.B2(n_1664),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1730),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1752),
.B(n_1705),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1718),
.B(n_1687),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1720),
.B(n_1692),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1719),
.B(n_1692),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1736),
.B(n_1571),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1737),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1724),
.B(n_1715),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1752),
.B(n_1637),
.C(n_1669),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1734),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1730),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1737),
.Y(n_1796)
);

NOR2x1p5_ASAP7_75t_L g1797 ( 
.A(n_1724),
.B(n_1565),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1717),
.A2(n_1697),
.B1(n_1672),
.B2(n_1669),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1758),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1756),
.B(n_1675),
.C(n_1717),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

CKINVDCx16_ASAP7_75t_R g1802 ( 
.A(n_1790),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1765),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1765),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1778),
.A2(n_1744),
.B1(n_1720),
.B2(n_1721),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1762),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1782),
.B(n_1719),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1784),
.B(n_1744),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1761),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1768),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1766),
.A2(n_1757),
.B(n_1786),
.C(n_1773),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1763),
.B(n_1721),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1775),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1768),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1763),
.Y(n_1815)
);

OAI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1798),
.A2(n_1686),
.B1(n_1748),
.B2(n_1750),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1764),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1764),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1782),
.B(n_1727),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1769),
.B(n_1729),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1727),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1761),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1794),
.B(n_1729),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1779),
.Y(n_1824)
);

OR2x6_ASAP7_75t_L g1825 ( 
.A(n_1770),
.B(n_1541),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1793),
.B(n_1744),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1779),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1769),
.B(n_1733),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1757),
.A2(n_1774),
.B1(n_1797),
.B2(n_1776),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1759),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1772),
.B(n_1733),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1781),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1781),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1759),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1799),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1818),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1800),
.A2(n_1826),
.B1(n_1815),
.B2(n_1808),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1811),
.A2(n_1770),
.B1(n_1783),
.B2(n_1787),
.C(n_1786),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1815),
.A2(n_1771),
.B1(n_1760),
.B2(n_1772),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1812),
.B(n_1760),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1806),
.B(n_1780),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1812),
.B(n_1773),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1792),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1799),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1803),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1817),
.A2(n_1792),
.B1(n_1777),
.B2(n_1795),
.C(n_1785),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1803),
.Y(n_1847)
);

OAI322xp33_ASAP7_75t_L g1848 ( 
.A1(n_1805),
.A2(n_1789),
.A3(n_1788),
.B1(n_1796),
.B2(n_1791),
.C1(n_1767),
.C2(n_1775),
.Y(n_1848)
);

OAI211xp5_ASAP7_75t_L g1849 ( 
.A1(n_1818),
.A2(n_1775),
.B(n_1501),
.C(n_1791),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1801),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1802),
.B(n_1792),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1809),
.B(n_1754),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1820),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1804),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1820),
.B(n_1754),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1828),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1822),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1829),
.A2(n_1686),
.B1(n_1789),
.B2(n_1723),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1828),
.B(n_1767),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1810),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1851),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1857),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1851),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1849),
.B(n_1841),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1843),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1840),
.B(n_1831),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1836),
.B(n_1837),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1857),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1840),
.B(n_1822),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1842),
.B(n_1831),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1843),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1860),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1853),
.B(n_1814),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1852),
.B(n_1807),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1853),
.B(n_1824),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1842),
.B(n_1825),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1860),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1835),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1856),
.Y(n_1879)
);

AND2x2_ASAP7_75t_SL g1880 ( 
.A(n_1846),
.B(n_1807),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1861),
.A2(n_1838),
.B(n_1839),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1865),
.B(n_1856),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1848),
.C(n_1850),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1879),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1880),
.B(n_1816),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1864),
.A2(n_1854),
.B(n_1847),
.C(n_1844),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1855),
.B1(n_1825),
.B2(n_1823),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1863),
.A2(n_1858),
.B1(n_1845),
.B2(n_1859),
.C(n_1832),
.Y(n_1888)
);

OA22x2_ASAP7_75t_L g1889 ( 
.A1(n_1865),
.A2(n_1825),
.B1(n_1813),
.B2(n_1859),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1871),
.A2(n_1827),
.B(n_1832),
.C(n_1810),
.Y(n_1890)
);

NAND4xp25_ASAP7_75t_L g1891 ( 
.A(n_1869),
.B(n_1833),
.C(n_1834),
.D(n_1830),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1870),
.B(n_1819),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1870),
.A2(n_1825),
.B(n_1833),
.Y(n_1893)
);

NAND4xp25_ASAP7_75t_L g1894 ( 
.A(n_1876),
.B(n_1834),
.C(n_1830),
.D(n_1819),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1884),
.B(n_1862),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1887),
.B(n_1866),
.Y(n_1896)
);

NAND4xp75_ASAP7_75t_L g1897 ( 
.A(n_1885),
.B(n_1868),
.C(n_1876),
.D(n_1866),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1882),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1881),
.B(n_1874),
.Y(n_1899)
);

NAND4xp25_ASAP7_75t_L g1900 ( 
.A(n_1883),
.B(n_1873),
.C(n_1875),
.D(n_1874),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1892),
.Y(n_1901)
);

OAI22xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1893),
.A2(n_1868),
.B1(n_1878),
.B2(n_1872),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1886),
.A2(n_1877),
.B(n_1872),
.C(n_1821),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1890),
.Y(n_1904)
);

NOR3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1894),
.B(n_1877),
.C(n_1492),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_SL g1906 ( 
.A(n_1899),
.B(n_1888),
.C(n_1492),
.Y(n_1906)
);

NAND3xp33_ASAP7_75t_SL g1907 ( 
.A(n_1904),
.B(n_1389),
.C(n_1889),
.Y(n_1907)
);

AOI21xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1896),
.A2(n_1821),
.B(n_1420),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1901),
.B(n_1501),
.C(n_1891),
.Y(n_1909)
);

NOR2xp67_ASAP7_75t_L g1910 ( 
.A(n_1900),
.B(n_1796),
.Y(n_1910)
);

AOI211xp5_ASAP7_75t_L g1911 ( 
.A1(n_1902),
.A2(n_1450),
.B(n_1694),
.C(n_1704),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1906),
.B(n_1897),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1910),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1908),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1909),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1907),
.A2(n_1898),
.B1(n_1905),
.B2(n_1895),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1910),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1912),
.B(n_1903),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_L g1921 ( 
.A(n_1915),
.B(n_1450),
.C(n_1477),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1912),
.B(n_1445),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1913),
.B(n_1918),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1917),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1919),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1922),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1923),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1925),
.Y(n_1928)
);

OAI211xp5_ASAP7_75t_SL g1929 ( 
.A1(n_1928),
.A2(n_1924),
.B(n_1916),
.C(n_1927),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1921),
.B1(n_1920),
.B2(n_1926),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1929),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1930),
.A2(n_1564),
.B(n_1477),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1931),
.A2(n_1743),
.B1(n_1732),
.B2(n_1704),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1932),
.A2(n_1743),
.B(n_1732),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1933),
.A2(n_1696),
.B(n_1694),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1934),
.A2(n_1536),
.B(n_1564),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_SL g1937 ( 
.A1(n_1936),
.A2(n_1935),
.B1(n_1536),
.B2(n_1570),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1704),
.B1(n_1694),
.B2(n_1702),
.C(n_1696),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1938),
.A2(n_1569),
.B(n_1570),
.C(n_1536),
.Y(n_1939)
);


endmodule