module fake_jpeg_49_n_596 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_596);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_596;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_57),
.B(n_97),
.Y(n_161)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_59),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_68),
.Y(n_124)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_1),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx2_ASAP7_75t_SL g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_96),
.Y(n_142)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_19),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_101),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_105),
.Y(n_168)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_30),
.B(n_47),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_28),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_43),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_51),
.B1(n_48),
.B2(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_112),
.A2(n_126),
.B1(n_138),
.B2(n_149),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_51),
.B1(n_48),
.B2(n_38),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_43),
.B1(n_54),
.B2(n_52),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_133),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_28),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_143),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_56),
.A2(n_37),
.B1(n_48),
.B2(n_31),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_145),
.B1(n_154),
.B2(n_157),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_47),
.B1(n_30),
.B2(n_38),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_136),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_22),
.B1(n_31),
.B2(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_41),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_71),
.A2(n_22),
.B1(n_37),
.B2(n_31),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_60),
.A2(n_51),
.B1(n_22),
.B2(n_54),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_84),
.A2(n_54),
.B1(n_52),
.B2(n_50),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_150),
.A2(n_160),
.B1(n_170),
.B2(n_172),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_43),
.C(n_50),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_151),
.B(n_165),
.C(n_7),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_91),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_27),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_64),
.A2(n_46),
.B1(n_44),
.B2(n_27),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_43),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_73),
.A2(n_44),
.B1(n_27),
.B2(n_41),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_175),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_75),
.B(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_93),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_76),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_76),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_78),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_58),
.A2(n_28),
.B1(n_43),
.B2(n_3),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_238)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_96),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_179),
.B(n_185),
.Y(n_283)
);

OR2x4_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_123),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_180),
.Y(n_273)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_181),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_182),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_183),
.B(n_184),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_109),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_123),
.A2(n_106),
.B1(n_100),
.B2(n_98),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_188),
.A2(n_164),
.B1(n_146),
.B2(n_171),
.Y(n_296)
);

OR2x4_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_43),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_189),
.A2(n_215),
.B(n_217),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_115),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_211),
.Y(n_263)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_240),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_196),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_92),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_203),
.Y(n_244)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_1),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_143),
.B(n_88),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_1),
.Y(n_210)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_2),
.C(n_3),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_226),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_133),
.A2(n_2),
.B(n_4),
.C(n_6),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_234),
.B(n_167),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_4),
.B(n_6),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g217 ( 
.A(n_138),
.B(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_152),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_116),
.A2(n_83),
.B1(n_81),
.B2(n_9),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_231),
.B1(n_159),
.B2(n_119),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_223),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_156),
.C(n_144),
.Y(n_243)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_132),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_7),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_229),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_114),
.B(n_8),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_118),
.B(n_144),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_235),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_129),
.A2(n_8),
.B(n_9),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_239),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_215),
.B1(n_234),
.B2(n_187),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_167),
.B1(n_146),
.B2(n_163),
.Y(n_274)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_113),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_241),
.A2(n_220),
.B1(n_177),
.B2(n_231),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_246),
.C(n_181),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_156),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_167),
.B1(n_140),
.B2(n_154),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_247),
.A2(n_17),
.B(n_19),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_116),
.B1(n_114),
.B2(n_174),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_288),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_137),
.B1(n_129),
.B2(n_174),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

AOI22x1_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_216),
.B1(n_189),
.B2(n_186),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_175),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_279),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_175),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_175),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_280),
.A2(n_266),
.B(n_285),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_194),
.A2(n_162),
.B1(n_153),
.B2(n_139),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_281),
.A2(n_17),
.B1(n_19),
.B2(n_263),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_188),
.B(n_162),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_285),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_125),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_137),
.B1(n_164),
.B2(n_163),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_225),
.B1(n_211),
.B2(n_221),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_239),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_242),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_317),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_311),
.B1(n_321),
.B2(n_330),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_218),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_301),
.B(n_304),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_206),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_313),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_244),
.B(n_191),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_259),
.B(n_198),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_307),
.B(n_315),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_335),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_209),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_324),
.C(n_292),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_273),
.A2(n_190),
.B(n_196),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_316),
.B(n_263),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_207),
.B1(n_219),
.B2(n_223),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_236),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_235),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_327),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_272),
.B(n_204),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_280),
.B(n_276),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_282),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

AOI22x1_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_182),
.B1(n_193),
.B2(n_227),
.Y(n_323)
);

OA22x2_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_247),
.B1(n_251),
.B2(n_296),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_243),
.B(n_200),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_201),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_13),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_328),
.B(n_329),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_242),
.B(n_14),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_19),
.B1(n_15),
.B2(n_16),
.Y(n_330)
);

INVx11_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_249),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_261),
.B1(n_254),
.B2(n_289),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_282),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_342),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_256),
.B(n_16),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_337),
.A2(n_241),
.B1(n_263),
.B2(n_265),
.Y(n_356)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_339),
.A2(n_343),
.B(n_347),
.Y(n_365)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_256),
.B(n_17),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_291),
.B(n_261),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_345),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_260),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_254),
.Y(n_346)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_266),
.A2(n_260),
.B(n_262),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_354),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_355),
.B(n_362),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_356),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_303),
.A2(n_288),
.B1(n_287),
.B2(n_264),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_366),
.A2(n_381),
.B1(n_326),
.B2(n_341),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_370),
.C(n_377),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_294),
.C(n_245),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_314),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_322),
.A2(n_287),
.B(n_289),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_384),
.B(n_310),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_245),
.C(n_286),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_303),
.A2(n_264),
.B1(n_293),
.B2(n_275),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_286),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_388),
.C(n_392),
.Y(n_407)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_383),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_316),
.A2(n_257),
.B(n_290),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_320),
.A2(n_269),
.B1(n_275),
.B2(n_293),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_387),
.A2(n_336),
.B1(n_317),
.B2(n_334),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_309),
.B(n_248),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_248),
.C(n_250),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_302),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_301),
.C(n_347),
.Y(n_418)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_402),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_396),
.A2(n_403),
.B1(n_418),
.B2(n_355),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_361),
.B(n_332),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_423),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_401),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_352),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_332),
.B1(n_328),
.B2(n_320),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_404),
.B(n_419),
.Y(n_461)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_405),
.Y(n_443)
);

HAxp5_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_345),
.CON(n_409),
.SN(n_409)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_409),
.A2(n_410),
.B(n_367),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_307),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_422),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_332),
.C(n_344),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_421),
.C(n_424),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_416),
.Y(n_437)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_335),
.Y(n_416)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_312),
.A3(n_304),
.B1(n_327),
.B2(n_315),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_420),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_364),
.B(n_329),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_371),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_350),
.B(n_312),
.C(n_338),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_342),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_340),
.C(n_323),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_370),
.B(n_323),
.C(n_346),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_392),
.C(n_382),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_354),
.A2(n_333),
.B1(n_330),
.B2(n_321),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_406),
.B1(n_430),
.B2(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_376),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_428),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_339),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_363),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_359),
.B(n_385),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_250),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_432),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_466),
.B1(n_396),
.B2(n_427),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_447),
.C(n_454),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_365),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_448),
.Y(n_474)
);

XNOR2x1_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_384),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_446),
.B(n_452),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_375),
.C(n_390),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_356),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_355),
.B(n_363),
.C(n_331),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_457),
.B(n_459),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_379),
.Y(n_453)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_358),
.C(n_389),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_407),
.B(n_358),
.C(n_386),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_467),
.C(n_433),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_398),
.A2(n_391),
.B(n_383),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_400),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_400),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_SL g459 ( 
.A1(n_430),
.A2(n_355),
.B(n_379),
.C(n_357),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_460),
.A2(n_417),
.B1(n_409),
.B2(n_415),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_353),
.Y(n_463)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_463),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g464 ( 
.A(n_413),
.B(n_380),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_429),
.C(n_416),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_410),
.A2(n_351),
.B(n_373),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_468),
.B(n_457),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_426),
.A2(n_353),
.B1(n_373),
.B2(n_368),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_368),
.C(n_367),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_401),
.Y(n_470)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_470),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_471),
.A2(n_477),
.B1(n_487),
.B2(n_490),
.Y(n_500)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_473),
.Y(n_511)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_439),
.Y(n_475)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_475),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_414),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_494),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_441),
.A2(n_425),
.B1(n_424),
.B2(n_398),
.Y(n_477)
);

AOI21xp33_ASAP7_75t_L g521 ( 
.A1(n_478),
.A2(n_449),
.B(n_459),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_420),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_483),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g507 ( 
.A1(n_481),
.A2(n_452),
.B(n_468),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_461),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_482),
.B(n_484),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_325),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_408),
.C(n_397),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_492),
.C(n_442),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_456),
.B(n_411),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_491),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_451),
.A2(n_405),
.B1(n_395),
.B2(n_360),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_348),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_434),
.B(n_360),
.C(n_391),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_436),
.B(n_306),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_493),
.B(n_496),
.Y(n_522)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_451),
.A2(n_269),
.B1(n_270),
.B2(n_290),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_447),
.B(n_270),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_497),
.A2(n_435),
.B(n_449),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_467),
.B(n_438),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_448),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_502),
.B(n_507),
.Y(n_537)
);

BUFx12_ASAP7_75t_L g504 ( 
.A(n_493),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_504),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_505),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_446),
.Y(n_508)
);

MAJx2_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_474),
.C(n_486),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_434),
.C(n_444),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_515),
.C(n_519),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_475),
.A2(n_466),
.B1(n_437),
.B2(n_435),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_513),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_518),
.B(n_488),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_435),
.C(n_437),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_483),
.B(n_445),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_517),
.B(n_496),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_497),
.A2(n_449),
.B(n_459),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_455),
.C(n_459),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_488),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_476),
.B(n_472),
.Y(n_523)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_515),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_520),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_485),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_525),
.B(n_531),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_501),
.A2(n_472),
.B1(n_477),
.B2(n_473),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_526),
.A2(n_536),
.B1(n_532),
.B2(n_511),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_528),
.B(n_503),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_529),
.A2(n_514),
.B(n_518),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_495),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_474),
.C(n_486),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_533),
.B(n_534),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_522),
.C(n_519),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_533),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_506),
.B1(n_516),
.B2(n_511),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_523),
.Y(n_551)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_469),
.C(n_494),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_534),
.C(n_530),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_544),
.A2(n_552),
.B(n_554),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_550),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_549),
.A2(n_551),
.B(n_541),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_509),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_555),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_527),
.B(n_520),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_499),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_537),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_556),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_469),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_558),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_504),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_540),
.A2(n_529),
.B(n_536),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_559),
.A2(n_551),
.B(n_550),
.Y(n_566)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_564),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_566),
.B(n_573),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_524),
.C(n_542),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_568),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_556),
.A2(n_538),
.B1(n_539),
.B2(n_526),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_560),
.A2(n_538),
.B1(n_539),
.B2(n_504),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_569),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_547),
.B(n_553),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_570),
.B(n_572),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_559),
.A2(n_549),
.B(n_555),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_546),
.A2(n_544),
.B(n_558),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_567),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_575),
.A2(n_565),
.B(n_583),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_572),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_561),
.C(n_569),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_562),
.B(n_563),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_SL g587 ( 
.A(n_578),
.B(n_579),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_564),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_L g589 ( 
.A(n_584),
.B(n_588),
.C(n_582),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_580),
.B(n_565),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_571),
.C(n_586),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_586),
.Y(n_590)
);

NAND4xp25_ASAP7_75t_L g588 ( 
.A(n_576),
.B(n_582),
.C(n_581),
.D(n_579),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_589),
.B(n_591),
.C(n_586),
.Y(n_593)
);

FAx1_ASAP7_75t_SL g592 ( 
.A(n_590),
.B(n_587),
.CI(n_585),
.CON(n_592),
.SN(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_592),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_593),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_593),
.Y(n_596)
);


endmodule