module fake_jpeg_24610_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_46),
.B1(n_49),
.B2(n_54),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_20),
.B1(n_36),
.B2(n_26),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_12),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_22),
.B1(n_24),
.B2(n_23),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_23),
.B1(n_20),
.B2(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_33),
.B1(n_19),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_39),
.B1(n_54),
.B2(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_63),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_70),
.B1(n_48),
.B2(n_53),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_58),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_72),
.B1(n_48),
.B2(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_93),
.B1(n_95),
.B2(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_87),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_74),
.B1(n_70),
.B2(n_62),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_47),
.B(n_40),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_76),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_64),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_50),
.B1(n_45),
.B2(n_40),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_111),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_83),
.B(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_106),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_80),
.B(n_78),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_70),
.B1(n_68),
.B2(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_77),
.B1(n_93),
.B2(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_131),
.B(n_107),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_126),
.B1(n_138),
.B2(n_113),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_124),
.B(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_116),
.B(n_97),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_68),
.B1(n_77),
.B2(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_98),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_80),
.B1(n_110),
.B2(n_55),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_83),
.B(n_85),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_121),
.B1(n_126),
.B2(n_138),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_90),
.B(n_85),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_50),
.B(n_69),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_64),
.B1(n_90),
.B2(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_157),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_143),
.Y(n_173)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_79),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_128),
.B1(n_123),
.B2(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_131),
.C(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_151),
.C(n_115),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_135),
.B1(n_104),
.B2(n_71),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_98),
.C(n_108),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_160),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_96),
.B1(n_104),
.B2(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_126),
.B1(n_121),
.B2(n_124),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_64),
.B(n_73),
.C(n_38),
.D(n_31),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_115),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_28),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_130),
.C(n_117),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.C(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_118),
.C(n_123),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_175),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_174),
.A2(n_162),
.B1(n_141),
.B2(n_156),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_112),
.B1(n_79),
.B2(n_81),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_79),
.B1(n_42),
.B2(n_15),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_28),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_146),
.B(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_32),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_181),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_166),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_149),
.B(n_183),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_188),
.B(n_193),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_158),
.B1(n_147),
.B2(n_155),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_19),
.B1(n_15),
.B2(n_25),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_158),
.B(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_176),
.B1(n_150),
.B2(n_174),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_145),
.C(n_142),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_34),
.C(n_25),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_157),
.C(n_154),
.Y(n_202)
);

OAI322xp33_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_166),
.A3(n_180),
.B1(n_139),
.B2(n_169),
.C1(n_163),
.C2(n_177),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_204),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_206),
.A2(n_210),
.B1(n_186),
.B2(n_193),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_42),
.B1(n_26),
.B2(n_25),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_209),
.B1(n_211),
.B2(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_214),
.C(n_194),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_199),
.B1(n_188),
.B2(n_200),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_214)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_220),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_0),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_212),
.B1(n_217),
.B2(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_230),
.B1(n_220),
.B2(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_203),
.B1(n_194),
.B2(n_4),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_215),
.B(n_218),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_2),
.C(n_3),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_3),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_244),
.B(n_241),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_210),
.B1(n_217),
.B2(n_215),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_242),
.B1(n_8),
.B2(n_9),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_7),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_212),
.C(n_219),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.C(n_6),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_5),
.C(n_6),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_6),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_7),
.C(n_8),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_9),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_10),
.B(n_11),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_263),
.B(n_10),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_238),
.B1(n_240),
.B2(n_245),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_249),
.B(n_248),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_10),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_261),
.B(n_260),
.Y(n_270)
);

OAI31xp33_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_269),
.A3(n_259),
.B(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_10),
.Y(n_273)
);


endmodule