module fake_jpeg_14674_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_0),
.B(n_3),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_10),
.B(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_9),
.C(n_14),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_7),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_11),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.C(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_29),
.B(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_46),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_21),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B(n_43),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.C(n_4),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.C(n_5),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_6),
.B(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_50),
.B1(n_0),
.B2(n_3),
.Y(n_58)
);


endmodule