module fake_jpeg_14035_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_60),
.B(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_77),
.Y(n_124)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_65),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_87),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_82),
.Y(n_165)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_18),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_21),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_21),
.B(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_103),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_32),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_45),
.B1(n_46),
.B2(n_25),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_106),
.A2(n_107),
.B(n_159),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_45),
.B1(n_46),
.B2(n_25),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_51),
.B1(n_22),
.B2(n_42),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_113),
.A2(n_140),
.B1(n_106),
.B2(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_53),
.B(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_58),
.B(n_29),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_135),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_52),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_44),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_69),
.A2(n_42),
.B1(n_45),
.B2(n_52),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_28),
.Y(n_150)
);

OR2x2_ASAP7_75t_SL g151 ( 
.A(n_65),
.B(n_24),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_24),
.B(n_28),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_23),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_19),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_88),
.A2(n_45),
.B1(n_32),
.B2(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_76),
.B(n_52),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_20),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_171),
.B(n_199),
.Y(n_238)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_178),
.B(n_185),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_103),
.B1(n_102),
.B2(n_100),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_186),
.Y(n_265)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_79),
.B1(n_97),
.B2(n_96),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_67),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_91),
.B1(n_86),
.B2(n_81),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_113),
.A2(n_146),
.B1(n_134),
.B2(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_188),
.A2(n_193),
.B1(n_43),
.B2(n_164),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_131),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

AO22x1_ASAP7_75t_SL g192 ( 
.A1(n_134),
.A2(n_20),
.B1(n_43),
.B2(n_68),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_202),
.B1(n_43),
.B2(n_110),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_42),
.B1(n_19),
.B2(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_82),
.B1(n_71),
.B2(n_66),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_203),
.B1(n_211),
.B2(n_218),
.Y(n_230)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_144),
.B(n_30),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_221),
.Y(n_235)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_198),
.B(n_200),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_139),
.B(n_67),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_138),
.A2(n_35),
.B(n_30),
.C(n_44),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_204),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_150),
.A2(n_42),
.B1(n_44),
.B2(n_30),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_205),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_255)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_207),
.Y(n_268)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_109),
.B(n_101),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_160),
.C(n_165),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_35),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_217),
.Y(n_262)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_35),
.B(n_20),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_190),
.B(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_105),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_223),
.Y(n_250)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_232),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_132),
.B1(n_143),
.B2(n_145),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_249),
.B1(n_257),
.B2(n_263),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_174),
.C(n_184),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_236),
.C(n_240),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_130),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_111),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_0),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_119),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_258),
.C(n_221),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_188),
.A2(n_121),
.B1(n_137),
.B2(n_161),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_180),
.A2(n_121),
.B1(n_137),
.B2(n_161),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_163),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_110),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_264),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_192),
.A2(n_164),
.B1(n_158),
.B2(n_125),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_261),
.A2(n_39),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_196),
.B(n_23),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_208),
.A2(n_157),
.B1(n_32),
.B2(n_23),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g272 ( 
.A1(n_201),
.A2(n_32),
.A3(n_23),
.B1(n_68),
.B2(n_98),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_23),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_32),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_193),
.B1(n_225),
.B2(n_203),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_283),
.B1(n_286),
.B2(n_304),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_202),
.B1(n_211),
.B2(n_220),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_279),
.A2(n_305),
.B1(n_317),
.B2(n_319),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_303),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_218),
.B1(n_206),
.B2(n_176),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_213),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_284),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_214),
.B1(n_172),
.B2(n_191),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_187),
.B1(n_173),
.B2(n_169),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_288),
.B(n_275),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_224),
.C(n_32),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_294),
.C(n_302),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_268),
.Y(n_290)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_290),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_0),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_233),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_226),
.B(n_228),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_292),
.A2(n_230),
.B(n_270),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g293 ( 
.A1(n_244),
.A2(n_0),
.B(n_1),
.Y(n_293)
);

AO21x2_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_252),
.B(n_247),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_234),
.B(n_39),
.C(n_1),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_250),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_300),
.Y(n_357)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_296),
.A2(n_311),
.B(n_321),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_250),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_9),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_39),
.C(n_1),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_9),
.C(n_18),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_255),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_229),
.A2(n_257),
.B1(n_228),
.B2(n_240),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_260),
.B1(n_246),
.B2(n_274),
.Y(n_359)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_244),
.A2(n_39),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_308)
);

XOR2x2_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_260),
.Y(n_361)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_238),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_271),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_245),
.A2(n_15),
.B(n_9),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_314),
.B(n_310),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_262),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_239),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_253),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_253),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_232),
.C(n_264),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_254),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_244),
.A2(n_14),
.B1(n_4),
.B2(n_6),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_233),
.B1(n_247),
.B2(n_242),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_332),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_325),
.B(n_328),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_295),
.B(n_239),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_337),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_297),
.A2(n_252),
.B1(n_227),
.B2(n_271),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_331),
.A2(n_297),
.B1(n_316),
.B2(n_290),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_282),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_352),
.C(n_281),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_338),
.A2(n_354),
.B(n_359),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_345),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_342),
.A2(n_347),
.B1(n_348),
.B2(n_361),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_356),
.B1(n_358),
.B2(n_329),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_282),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_305),
.A2(n_267),
.B1(n_227),
.B2(n_231),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_248),
.B1(n_269),
.B2(n_256),
.Y(n_348)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_296),
.A3(n_288),
.B1(n_300),
.B2(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_351),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_299),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_248),
.Y(n_352)
);

A2O1A1O1Ixp25_ASAP7_75t_L g354 ( 
.A1(n_277),
.A2(n_292),
.B(n_280),
.C(n_320),
.D(n_285),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_276),
.A2(n_269),
.B1(n_251),
.B2(n_256),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_356),
.A2(n_358),
.B1(n_278),
.B2(n_279),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_283),
.A2(n_251),
.B1(n_241),
.B2(n_243),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_290),
.B(n_273),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_362),
.A2(n_353),
.B(n_338),
.Y(n_392)
);

OAI21x1_ASAP7_75t_R g364 ( 
.A1(n_344),
.A2(n_293),
.B(n_306),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_364),
.A2(n_367),
.B(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_324),
.A2(n_296),
.B1(n_304),
.B2(n_281),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_376),
.B1(n_383),
.B2(n_384),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_332),
.A2(n_293),
.B1(n_278),
.B2(n_294),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_380),
.B1(n_385),
.B2(n_395),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_381),
.C(n_393),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_281),
.B1(n_293),
.B2(n_309),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_357),
.A2(n_293),
.A3(n_318),
.B1(n_298),
.B2(n_303),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_388),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_289),
.B(n_274),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_345),
.A2(n_312),
.B1(n_302),
.B2(n_319),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_317),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_361),
.A2(n_347),
.B1(n_348),
.B2(n_342),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_315),
.B1(n_246),
.B2(n_273),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_360),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_337),
.B(n_3),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_387),
.Y(n_410)
);

AOI31xp33_ASAP7_75t_SL g388 ( 
.A1(n_349),
.A2(n_4),
.A3(n_6),
.B(n_7),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_330),
.A2(n_7),
.A3(n_328),
.B1(n_353),
.B2(n_343),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_391),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_360),
.A2(n_7),
.B1(n_355),
.B2(n_336),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_326),
.C(n_350),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_336),
.A2(n_322),
.B1(n_344),
.B2(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_323),
.B(n_339),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_396),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_344),
.B(n_339),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_397),
.A2(n_362),
.B(n_344),
.Y(n_406)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_405),
.Y(n_448)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_350),
.C(n_326),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_412),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_335),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_406),
.A2(n_397),
.B(n_392),
.Y(n_445)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_389),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_408),
.B(n_386),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_419),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_354),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_414),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_389),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_335),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_365),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_381),
.B(n_333),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_425),
.Y(n_432)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_374),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_374),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_333),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_378),
.C(n_414),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_455),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_399),
.A2(n_394),
.B1(n_372),
.B2(n_363),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_434),
.A2(n_437),
.B1(n_440),
.B2(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_363),
.B1(n_383),
.B2(n_391),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_398),
.A2(n_413),
.B1(n_417),
.B2(n_427),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_409),
.A2(n_395),
.B1(n_371),
.B2(n_366),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_445),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_425),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_413),
.A2(n_376),
.B1(n_368),
.B2(n_384),
.Y(n_443)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_380),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_447),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_411),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_409),
.A2(n_385),
.B1(n_377),
.B2(n_364),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_454),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_367),
.C(n_327),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_453),
.C(n_431),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_327),
.C(n_351),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_419),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_422),
.B(n_429),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_439),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_457),
.B(n_473),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_459),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_451),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_470),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g465 ( 
.A1(n_456),
.A2(n_454),
.B(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_403),
.C(n_421),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_469),
.C(n_477),
.Y(n_481)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_430),
.C(n_432),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_443),
.A2(n_421),
.B1(n_398),
.B2(n_417),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_472),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_426),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_426),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_L g475 ( 
.A1(n_445),
.A2(n_424),
.B(n_404),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_475),
.A2(n_452),
.B(n_404),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_401),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_390),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_401),
.C(n_406),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_475),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_441),
.C(n_434),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_484),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_437),
.C(n_435),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_435),
.C(n_433),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_487),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_433),
.C(n_449),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_461),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_491),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_344),
.B1(n_407),
.B2(n_450),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_462),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_460),
.A2(n_450),
.B(n_438),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_490),
.A2(n_410),
.B1(n_423),
.B2(n_420),
.Y(n_509)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_463),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_474),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_484),
.C(n_487),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_501),
.Y(n_515)
);

OR2x6_ASAP7_75t_SL g514 ( 
.A(n_498),
.B(n_480),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_472),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_509),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_458),
.C(n_477),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_503),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_444),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_504),
.B(n_507),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_467),
.C(n_470),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_510),
.C(n_501),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_467),
.C(n_438),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_485),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_493),
.C(n_492),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_505),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_512),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_506),
.A2(n_483),
.B1(n_494),
.B2(n_490),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_483),
.B1(n_465),
.B2(n_415),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_514),
.Y(n_525)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_522),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_498),
.A2(n_410),
.B(n_388),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_388),
.B(n_364),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_341),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_517),
.A2(n_510),
.B(n_500),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_SL g530 ( 
.A1(n_526),
.A2(n_515),
.B(n_519),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_529),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_499),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_529),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_525),
.A2(n_512),
.B(n_516),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_531),
.A2(n_532),
.B(n_514),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_523),
.A2(n_514),
.B(n_521),
.Y(n_532)
);

AOI21x1_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_524),
.B(n_527),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_534),
.A2(n_536),
.B(n_520),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_535),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_537),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_538),
.C(n_528),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_400),
.C(n_340),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_364),
.Y(n_542)
);


endmodule