module fake_jpeg_1311_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_49),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_48),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_15),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_22),
.B1(n_33),
.B2(n_26),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_18),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_21),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_44),
.B1(n_39),
.B2(n_2),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_70),
.B1(n_45),
.B2(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_44),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_17),
.Y(n_70)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_8),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_88),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_45),
.B(n_34),
.C(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_34),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_55),
.B1(n_39),
.B2(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_12),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_58),
.B1(n_71),
.B2(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_77),
.B1(n_98),
.B2(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_112),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_52),
.A3(n_44),
.B1(n_39),
.B2(n_72),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_64),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_85),
.C(n_99),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_127),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_132),
.B1(n_135),
.B2(n_115),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_130),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_90),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_83),
.B1(n_94),
.B2(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_78),
.B1(n_93),
.B2(n_55),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_101),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_103),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_64),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_117),
.C(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_134),
.B1(n_132),
.B2(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_136),
.C(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_135),
.C(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_113),
.B(n_106),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_119),
.C(n_117),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_126),
.C(n_108),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_147),
.C(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_161),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_111),
.B1(n_104),
.B2(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_105),
.B1(n_102),
.B2(n_2),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_163),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_170),
.C(n_171),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_143),
.B(n_151),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_138),
.C(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_105),
.C(n_141),
.Y(n_171)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_154),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.C(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_0),
.C(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_165),
.Y(n_180)
);

OAI221xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_168),
.B1(n_102),
.B2(n_3),
.C(n_4),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_176),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_177),
.B(n_4),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_5),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_187),
.B(n_184),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_5),
.Y(n_190)
);


endmodule