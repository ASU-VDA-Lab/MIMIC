module fake_jpeg_21874_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_43),
.Y(n_66)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_57),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_33),
.B1(n_23),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_18),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_23),
.C(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_27),
.Y(n_95)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_33),
.B1(n_18),
.B2(n_21),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_33),
.B1(n_21),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_80),
.B1(n_88),
.B2(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_27),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_32),
.B(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_33),
.B1(n_26),
.B2(n_34),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_21),
.B1(n_26),
.B2(n_30),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_20),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_17),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_65),
.B1(n_48),
.B2(n_17),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_97),
.B(n_89),
.Y(n_151)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_120),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_11),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_102),
.C(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_45),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_57),
.C(n_49),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_10),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_111),
.B(n_74),
.Y(n_127)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_67),
.B1(n_51),
.B2(n_50),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_80),
.B1(n_71),
.B2(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_80),
.Y(n_128)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_48),
.B1(n_60),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_70),
.A2(n_48),
.B1(n_32),
.B2(n_17),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_27),
.C(n_20),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_72),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_131),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_129),
.B(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_103),
.B1(n_120),
.B2(n_107),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_141),
.B1(n_148),
.B2(n_86),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_91),
.B(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_145),
.B(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_149),
.B1(n_152),
.B2(n_82),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_92),
.B(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_88),
.B1(n_73),
.B2(n_96),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_73),
.B1(n_76),
.B2(n_86),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_106),
.C(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_158),
.C(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_124),
.C(n_118),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_116),
.B1(n_111),
.B2(n_97),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_164),
.B(n_167),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_182),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_112),
.B(n_114),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_173),
.B(n_181),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_112),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_76),
.B(n_94),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_145),
.C(n_132),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_175),
.C(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_121),
.C(n_69),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_86),
.B1(n_79),
.B2(n_82),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_185),
.B1(n_149),
.B2(n_129),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_99),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_109),
.B(n_69),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_184),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_147),
.C(n_150),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_168),
.C(n_165),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_133),
.C(n_126),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_208),
.B(n_11),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_204),
.B1(n_184),
.B2(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_141),
.B1(n_136),
.B2(n_134),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_177),
.B1(n_185),
.B2(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_134),
.C(n_135),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_190),
.C(n_191),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_130),
.B1(n_131),
.B2(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_209),
.Y(n_213)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_11),
.B(n_16),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_159),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_225),
.B1(n_232),
.B2(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_172),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_219),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_221),
.B(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_235),
.C(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_179),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_180),
.B(n_156),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_169),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_175),
.B1(n_167),
.B2(n_161),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_28),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_28),
.C(n_25),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_250),
.Y(n_267)
);

AOI321xp33_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_196),
.A3(n_194),
.B1(n_199),
.B2(n_200),
.C(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_220),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_194),
.C(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_245),
.C(n_249),
.Y(n_269)
);

AOI221xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_210),
.B1(n_188),
.B2(n_193),
.C(n_212),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_247),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_217),
.C(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_202),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_195),
.C(n_202),
.Y(n_249)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_257),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_195),
.C(n_187),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_229),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_265),
.C(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_234),
.B1(n_226),
.B2(n_233),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_270),
.B1(n_0),
.B2(n_1),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_223),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_9),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_256),
.B(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_213),
.B(n_226),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_252),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_228),
.Y(n_273)
);

OAI321xp33_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_22),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C(n_12),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_240),
.Y(n_274)
);

FAx1_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_254),
.CI(n_243),
.CON(n_276),
.SN(n_276)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_274),
.B(n_15),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_238),
.B1(n_245),
.B2(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_238),
.C(n_239),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_265),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_250),
.B1(n_232),
.B2(n_206),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_252),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_212),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_287),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_285),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_9),
.B(n_16),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_10),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_22),
.B(n_1),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_269),
.B(n_271),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_272),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_300),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_284),
.B1(n_285),
.B2(n_276),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_0),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_307),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_309),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_276),
.B(n_277),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_291),
.A3(n_275),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_5),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_297),
.B(n_293),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_315),
.B(n_4),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_312),
.A3(n_306),
.B1(n_5),
.B2(n_6),
.C1(n_4),
.C2(n_305),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_275),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_5),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_2),
.B(n_4),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_313),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_317),
.B(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_4),
.Y(n_321)
);


endmodule