module fake_jpeg_18963_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_32),
.B1(n_40),
.B2(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_28),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_48),
.B(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_50),
.B1(n_30),
.B2(n_24),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_77),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_15),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_41),
.B1(n_34),
.B2(n_18),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_72),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_16),
.B1(n_30),
.B2(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_19),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_36),
.B1(n_35),
.B2(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_39),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_35),
.B1(n_24),
.B2(n_15),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_10),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_48),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_55),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_14),
.B(n_13),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_48),
.B1(n_46),
.B2(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_54),
.C(n_25),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_90),
.C(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_108),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_83),
.B(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_111),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_15),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_67),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_73),
.B(n_68),
.C(n_58),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_89),
.B1(n_82),
.B2(n_67),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_27),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_15),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_91),
.C(n_81),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_83),
.B1(n_85),
.B2(n_81),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_138),
.B1(n_140),
.B2(n_107),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_111),
.C(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_113),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_139),
.B(n_29),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_89),
.B(n_15),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_126),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_155),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_116),
.B1(n_109),
.B2(n_123),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_113),
.A3(n_105),
.B1(n_108),
.B2(n_122),
.C1(n_29),
.C2(n_21),
.Y(n_149)
);

OAI322xp33_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_159),
.A3(n_21),
.B1(n_157),
.B2(n_156),
.C1(n_143),
.C2(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_157),
.B(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_133),
.B1(n_141),
.B2(n_129),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_29),
.B1(n_21),
.B2(n_5),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_2),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_8),
.C(n_14),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_166),
.Y(n_178)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_135),
.C(n_134),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_146),
.C(n_168),
.Y(n_172)
);

XOR2x2_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_144),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_151),
.B(n_144),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_153),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_3),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_179),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_162),
.B(n_6),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_163),
.C(n_169),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_177),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_9),
.C(n_11),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_3),
.C(n_5),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_185),
.B(n_5),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_162),
.B1(n_164),
.B2(n_7),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_187),
.Y(n_190)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_176),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_189),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_187),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_184),
.C(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_7),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_196),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_191),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_194),
.Y(n_199)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_200),
.B(n_190),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_202),
.Y(n_203)
);


endmodule