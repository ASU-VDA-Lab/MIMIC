module fake_jpeg_1419_n_75 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_43),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_32),
.B1(n_22),
.B2(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_22),
.C(n_20),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_38),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_51),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_38),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_R g53 ( 
.A(n_42),
.B(n_19),
.Y(n_53)
);

XNOR2x1_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_56),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_3),
.B(n_4),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_59),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_11),
.C(n_6),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_66),
.B1(n_64),
.B2(n_10),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_8),
.B(n_9),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_9),
.Y(n_75)
);


endmodule