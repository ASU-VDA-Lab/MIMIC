module fake_jpeg_490_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2x1_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_0),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.CON(n_91),
.SN(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_66),
.Y(n_89)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_71),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_65),
.B1(n_76),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_96),
.B1(n_79),
.B2(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_77),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_65),
.B1(n_76),
.B2(n_54),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_79),
.B1(n_84),
.B2(n_83),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_113),
.Y(n_119)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_81),
.B1(n_80),
.B2(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_110),
.B1(n_112),
.B2(n_103),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_81),
.B1(n_69),
.B2(n_60),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_85),
.B1(n_98),
.B2(n_59),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_26),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_60),
.B1(n_57),
.B2(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_57),
.B1(n_75),
.B2(n_56),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_56),
.B(n_53),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_64),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_67),
.C(n_55),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_62),
.C(n_5),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_133),
.B1(n_134),
.B2(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_73),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_8),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_95),
.B1(n_58),
.B2(n_61),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_61),
.B1(n_95),
.B2(n_62),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_144),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_62),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_42),
.C(n_41),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_95),
.B1(n_5),
.B2(n_6),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_155),
.B1(n_156),
.B2(n_18),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_154),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_52),
.B1(n_50),
.B2(n_49),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_4),
.B(n_6),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_139),
.B(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_11),
.B(n_12),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_162),
.B(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_11),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_13),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_163),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_14),
.B(n_15),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_176),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_137),
.B(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_148),
.A3(n_143),
.B1(n_156),
.B2(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_162),
.B1(n_152),
.B2(n_158),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_173),
.B1(n_168),
.B2(n_166),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_34),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_164),
.C(n_159),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_173),
.B1(n_181),
.B2(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_179),
.B1(n_169),
.B2(n_167),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_176),
.B1(n_152),
.B2(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_200),
.C(n_184),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_185),
.C(n_171),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_189),
.C(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_32),
.C(n_31),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_30),
.B(n_29),
.C(n_28),
.Y(n_206)
);

NAND4xp25_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_208),
.C(n_18),
.D(n_20),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_195),
.B1(n_19),
.B2(n_20),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_207),
.B(n_22),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_21),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_24),
.B(n_21),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_23),
.B(n_24),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_23),
.Y(n_215)
);


endmodule